----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:06:27 01/19/2019 
-- Design Name: 
-- Module Name:    ControlLogic - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ControlLogic is
    Port ( CLK : in STD_LOGIC;
           nRST : in STD_LOGIC;
           IReg : in STD_LOGIC_VECTOR (15 downto 0);
           ACval, DRval : in STD_LOGIC_VECTOR (15 downto 0);
           Eval : in STD_LOGIC;
           FGItoCL, FGOtoCL : in STD_LOGIC;
           FGInRST, FGOnRST : out STD_LOGIC;
           ArbiterSEL : out STD_LOGIC_VECTOR (2 downto 0);
           ARnRST, PCnRST, DRnRST, EnRST, ACnRST, INPRnRST, IRnRST, RegBanknRST, OUTRnRST : out STD_LOGIC;
           ARLD, PCLD, DRLD, ACLD, INPRLD, IRLD, OUTRLD : out STD_LOGIC;
           ARInc, PCInc, DRInc, ACInc, INPRInc, IRInc, OUTRInc : out STD_LOGIC;
           Ecmpl, ACcmpl : out STD_LOGIC;
           ALUfunc : out STD_LOGIC_VECTOR (3 downto 0);
           DRMUXSel, ACMUXSel : out STD_LOGIC;
           MemWR, MemRE : out STD_LOGIC;
           RegBankaddr : out STD_LOGIC_VECTOR (2 downto 0);
           RegBankRW : out STD_LOGIC;
           RegBankImmVal : out STD_LOGIC_VECTOR (7 downto 0);
           RegBankImmEn : out STD_LOGIC);
end ControlLogic;

architecture Behavioral of ControlLogic is

    type state is (T0, T1, T2, T3, T4, T5, T6, T7);
    signal pr_state, nx_state : state;

    signal ArbiterSELt : STD_LOGIC_VECTOR (2 downto 0) := "000";
    signal ARnRSTt, PCnRSTt, DRnRSTt, EnRSTt, ACnRSTt, INPRnRSTt, IRnRSTt, RegBanknRSTt, OUTRnRSTt : STD_LOGIC := '0';
    signal ARLDt, PCLDt, DRLDt, ACLDt, INPRLDt, IRLDt, OUTRLDt : STD_LOGIC := '0';
    signal ARInct, PCInct, DRInct, ACInct, INPRInct, IRInct, OUTRInct : STD_LOGIC := '0';
    signal Ecmplt, ACcmplt : STD_LOGIC := '0';
    signal ALUfunct : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal DRMUXSelt, ACMUXSelt : STD_LOGIC := '0';
    signal MemWRt, MemREt : STD_LOGIC := '0';
    signal RegBankaddrt : STD_LOGIC_VECTOR (2 downto 0) := "000";
    signal RegBankRWt : STD_LOGIC := '0';
    signal RegBankImmValt : STD_LOGIC_VECTOR (7 downto 0) := "00000000";
    signal RegBankImmEnt : STD_LOGIC := '0';

    signal memInstOpcode, ImmInstOpcode : STD_LOGIC_VECTOR (2 downto 0) := "000";
    signal RegInstOpcode : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal FGInRSTt, FGOnRSTt : STD_LOGIC := '1';
    signal RInt : STD_LOGIC := '0';

begin

    process (CLK, nRST)
    begin
        if (nRST = '0') then
            pr_state <= T0;
        elsif (rising_edge(CLK)) then
            pr_state <= nx_state;
        end if;
    end process;

    process (pr_state, IReg, ACval, DRval, Eval, FGItoCL, FGOtoCL)
    begin
        case (pr_state) is
            when T0 =>
                if (RInt = '1') then
                    ArbiterSELt <= "100"; --changed
                    ARnRSTt <= '1';
                    PCnRSTt <= '1';
                    DRnRSTt <= '1';
                    EnRSTt <= '1';
                    ACnRSTt <= '1';
                    INPRnRSTt <= '1';
                    IRnRSTt <= '1';
                    RegBanknRSTt <= '1';
                    OUTRnRSTt <= '1';
                    ARLDt <= '0';
                    PCLDt <= '0';
                    DRLDt <= '0';
                    ACLDt <= '0';
                    INPRLDt <= '0';
                    IRLDt <= '0';
                    OUTRLDt <= '0';
                    ARInct <= '0';
                    PCInct <= '0';
                    DRInct <= '0';
                    ACInct <= '0';
                    INPRInct <= '0';
                    IRInct <= '0';
                    OUTRInct <= '0';
                    Ecmplt <= '0';
                    ACcmplt <= '0';
                    ALUfunct <= "0000";
                    DRMUXSelt <= '0';
                    ACMUXSelt <= '0';
                    MemWRt <= '0';
                    MemREt <= '0';
                    RegBankaddrt <= "000"; --changed
                    RegBankRWt <= '1'; --changed
                    RegBankImmValt <= "00000000";
                    RegBankImmEnt <= '0';
                    FGInRSTt <= '1';
                    FGOnRSTt <= '1';
                    nx_state <= T1;
                else
                    ArbiterSELt <= "100"; --changed
                    ARnRSTt <= '1';
                    PCnRSTt <= '1';
                    DRnRSTt <= '1';
                    EnRSTt <= '1';
                    ACnRSTt <= '1';
                    INPRnRSTt <= '1';
                    IRnRSTt <= '1';
                    RegBanknRSTt <= '1';
                    OUTRnRSTt <= '1';
                    ARLDt <= '1'; --changed
                    PCLDt <= '0';
                    DRLDt <= '0';
                    ACLDt <= '0';
                    INPRLDt <= '0';
                    IRLDt <= '0';
                    OUTRLDt <= '0';
                    ARInct <= '0';
                    PCInct <= '0';
                    DRInct <= '0';
                    ACInct <= '0';
                    INPRInct <= '0';
                    IRInct <= '0';
                    OUTRInct <= '0';
                    Ecmplt <= '0';
                    ACcmplt <= '0';
                    ALUfunct <= "0000";
                    DRMUXSelt <= '0';
                    ACMUXSelt <= '0';
                    MemWRt <= '0';
                    MemREt <= '0';
                    RegBankaddrt <= "000";
                    RegBankRWt <= '0';
                    RegBankImmValt <= "00000000";
                    RegBankImmEnt <= '0';
                    FGInRSTt <= '1';
                    FGOnRSTt <= '1';
                    nx_state <= T1;
                end if;
            when T1 =>
                if (RInt = '1') then
                    RInt <= '0'; --changed
                    ArbiterSELt <= "000";
                    ARnRSTt <= '1';
                    PCnRSTt <= '0'; --changed
                    DRnRSTt <= '1';
                    EnRSTt <= '1';
                    ACnRSTt <= '1';
                    INPRnRSTt <= '1';
                    IRnRSTt <= '1';
                    RegBanknRSTt <= '1';
                    OUTRnRSTt <= '1';
                    ARLDt <= '0';
                    PCLDt <= '0';
                    DRLDt <= '0';
                    ACLDt <= '0';
                    INPRLDt <= '0';
                    IRLDt <= '0';
                    OUTRLDt <= '0';
                    ARInct <= '0';
                    PCInct <= '0';
                    DRInct <= '0';
                    ACInct <= '0';
                    INPRInct <= '0';
                    IRInct <= '0';
                    OUTRInct <= '0';
                    Ecmplt <= '0';
                    ACcmplt <= '0';
                    ALUfunct <= "0000";
                    DRMUXSelt <= '0';
                    ACMUXSelt <= '0';
                    MemWRt <= '0';
                    MemREt <= '0';
                    RegBankaddrt <= "000";
                    RegBankRWt <= '0';
                    RegBankImmValt <= "00000000";
                    RegBankImmEnt <= '0';
                    FGInRSTt <= '1';
                    FGOnRSTt <= '1';
                    nx_state <= T0;
                else
                    ArbiterSELt <= "110"; --changed
                    ARnRSTt <= '1';
                    PCnRSTt <= '1';
                    DRnRSTt <= '1';
                    EnRSTt <= '1';
                    ACnRSTt <= '1';
                    INPRnRSTt <= '1';
                    IRnRSTt <= '1';
                    RegBanknRSTt <= '1';
                    OUTRnRSTt <= '1';
                    ARLDt <= '0';
                    PCLDt <= '0';
                    DRLDt <= '0';
                    ACLDt <= '0';
                    INPRLDt <= '0';
                    IRLDt <= '1'; --changed
                    OUTRLDt <= '0';
                    ARInct <= '0';
                    PCInct <= '1'; --changed
                    DRInct <= '0';
                    ACInct <= '0';
                    INPRInct <= '0';
                    IRInct <= '0';
                    OUTRInct <= '0';
                    Ecmplt <= '0';
                    ACcmplt <= '0';
                    ALUfunct <= "0000";
                    DRMUXSelt <= '0';
                    ACMUXSelt <= '0';
                    MemWRt <= '0';
                    MemREt <= '1'; --changed
                    RegBankaddrt <= "000";
                    RegBankRWt <= '0';
                    RegBankImmValt <= "00000000";
                    RegBankImmEnt <= '0';
                    FGInRSTt <= '1';
                    FGOnRSTt <= '1';
                    nx_state <= T2;
                end if;
            when T2 =>
                if (FGItoCL = '1' or FGOtoCL = '1') then
                    RInt <= '1';
                else
                    RInt <= '0';
                end if;
                if (IReg(15) = '0') then -- memory instruction
                    memInstOpcode <= IReg(14 downto 12);
                else
                    if (IReg(14) = '0') then -- register instruction
                        RegInstOpcode <= IReg(13 downto 10);
                    else -- immediate instruction
                        ImmInstOpcode <= IReg(13 downto 11);
                    end if;
                end if;
                ArbiterSELt <= "010"; --changed
                ARnRSTt <= '1';
                PCnRSTt <= '1';
                DRnRSTt <= '1';
                EnRSTt <= '1';
                ACnRSTt <= '1';
                INPRnRSTt <= '1';
                IRnRSTt <= '1';
                RegBanknRSTt <= '1';
                OUTRnRSTt <= '1';
                ARLDt <= '1'; --changed
                PCLDt <= '0';
                DRLDt <= '0';
                ACLDt <= '0';
                INPRLDt <= '0';
                IRLDt <= '0';
                OUTRLDt <= '0';
                ARInct <= '0';
                PCInct <= '0';
                DRInct <= '0';
                ACInct <= '0';
                INPRInct <= '0';
                IRInct <= '0';
                OUTRInct <= '0';
                Ecmplt <= '0';
                ACcmplt <= '0';
                ALUfunct <= "0000";
                DRMUXSelt <= '0';
                ACMUXSelt <= '0';
                MemWRt <= '0';
                MemREt <= '0';
                RegBankaddrt <= "000";
                RegBankRWt <= '0';
                RegBankImmValt <= "00000000";
                RegBankImmEnt <= '0';
                FGInRSTt <= '1';
                FGOnRSTt <= '1';
                nx_state <= T3;
            when T3 =>
                if (IReg(15) = '0') then -- memory instruction
                    case (memInstOpcode) is
                        when "000" => -- ADD
                            ArbiterSELt <= "110"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '1'; --changed
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '1'; --changed
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when "001" => -- NAND
                            ArbiterSELt <= "110"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '1'; --changed
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '1'; --changed
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when "010" => -- NOT
                            ArbiterSELt <= "110"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '1'; --changed
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '1'; --changed
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when "011" => -- LDA
                            ArbiterSELt <= "110"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '1'; --changed
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '1'; --changed
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when "100" => -- STA
                            ArbiterSELt <= "001"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '1'; --changed
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "101" => -- BUN
                            ArbiterSELt <= "101"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '1'; --changed
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "110" => -- BSA
                            ArbiterSELt <= "100"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '1'; --changed
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '1'; --changed
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when "111" => -- ISZ
                            ArbiterSELt <= "110"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '1'; --changed
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '1'; --changed
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T4;
                        when others =>
                    end case;
                else
                    if (IReg(14) = '0') then -- register instruction
                        case (RegInstOpcode) is
                            when "0000" => -- ADDR
                                ArbiterSELt <= "011"; --changed
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '1'; --changed
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= IReg(6 downto 4); --changed
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T4;
                            when "0001" => -- SHR
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0100"; --changed
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '1'; --changed
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0010" => -- SHL
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0101"; --changed
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '1'; --changed
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0011" => -- CIR
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0110"; --changed
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '1'; --changed
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0100" => -- CIL
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0111"; --changed
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '1'; --changed
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0101" => -- INC
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '1'; --changed
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0110" => -- CLA
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '0'; --changed
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "0111" => -- CMA
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '1'; --changed
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1000" => -- CLE
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '0'; --changed
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1001" => -- CME
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '1'; --changed
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1010" => -- SZA
                                if (ACval = "0000000000000000") then
                                    PCInct <= '1'; --changed
                                else
                                    PCInct <= '0'; --changed
                                end if;
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1011" => -- SZE
                                if (Eval = '0') then
                                    PCInct <= '1'; --changed
                                else
                                    PCInct <= '0'; --changed
                                end if;
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1100" => -- INP
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "1000"; --changed
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '0'; --changed
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "1101" => -- OUT
                                ArbiterSELt <= "001"; --changed
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '1'; --changed
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= "000";
                                RegBankRWt <= '0';
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '0'; --changed
                                nx_state <= T0;
                            when others =>
                        end case;
                    else -- immediate instruction
                        case (ImmInstOpcode) is
                            when "000" => -- LDI
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= IReg(10 downto 8); --changed
                                RegBankRWt <= '1'; --changed
                                RegBankImmValt <= IReg(7 downto 0); --changed
                                RegBankImmEnt <= '1'; --changed
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when "001" => -- ADDI
                                ArbiterSELt <= "011"; --changed
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '1'; --changed
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= IReg(10 downto 8); --changed
                                RegBankRWt <= '0'; --changed
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T0;
                            when others =>
                        end case;
                    end if;
                end if;
            when T4 =>
                if (IReg(15) = '0') then -- memory instruction
                    case (memInstOpcode) is
                        when "000" => -- ADD
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '1'; --changed
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000"; --changed
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '1'; --changed
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "001" => -- NAND
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '1'; --changed
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0001"; --changed
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '1'; --changed
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "010" => -- NOT
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '1'; --changed
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "1001"; --changed
                            DRMUXSelt <= '0'; --changed
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "011" => -- LDA
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '1'; --changed
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0011"; --changed
                            DRMUXSelt <= '0'; --changed
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "110" => -- BSA
                            ArbiterSELt <= "101"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '1'; --changed
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when "111" => -- ISZ
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '1'; --changed
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T5;
                        when others =>
                    end case;
                else
                    if (IReg(14) = '0') then -- register instruction
                        case (RegInstOpcode) is
                            when "0000" => -- ADDR
                            ArbiterSELt <= "000";
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '1'; --changed
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000"; --changed
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '1'; --changed
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T5;
                            when others =>
                        end case;
                    else -- immediate instruction
                        case (ImmInstOpcode) is
                            when "001" => -- ADDI
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '0';
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000";
                                DRMUXSelt <= '0';
                                ACMUXSelt <= '0';
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= IReg(10 downto 8); --changed
                                RegBankRWt <= '1'; --changed
                                RegBankImmValt <= IReg(7 downto 0); --changed
                                RegBankImmEnt <= '1'; --changed
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T5;
                            when others =>
                        end case;
                    end if;
                end if;
            when T5 =>
                if (IReg(15) = '0') then -- memory instruction
                    case (memInstOpcode) is
                        when "111" => -- ISZ
                            if (DRval = "0000000000000000") then
                                PCInct <= '1'; --changed
                            else
                                PCInct <= '0'; --changed
                            end if;
                            ArbiterSELt <= "000"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '1'; --changed
                            MemREt <= '0';
                            RegBankaddrt <= "000";
                            RegBankRWt <= '0';
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                        when others =>
                    end case;
                else
                    if (IReg(14) = '0') then -- register instruction
                        case (RegInstOpcode) is
                            when "0000" => -- ADDR
                            ArbiterSELt <= "001"; --changed
                            ARnRSTt <= '1';
                            PCnRSTt <= '1';
                            DRnRSTt <= '1';
                            EnRSTt <= '1';
                            ACnRSTt <= '1';
                            INPRnRSTt <= '1';
                            IRnRSTt <= '1';
                            RegBanknRSTt <= '1';
                            OUTRnRSTt <= '1';
                            ARLDt <= '0';
                            PCLDt <= '0';
                            DRLDt <= '0';
                            ACLDt <= '0';
                            INPRLDt <= '0';
                            IRLDt <= '0';
                            OUTRLDt <= '0';
                            ARInct <= '0';
                            PCInct <= '0';
                            DRInct <= '0';
                            ACInct <= '0';
                            INPRInct <= '0';
                            IRInct <= '0';
                            OUTRInct <= '0';
                            Ecmplt <= '0';
                            ACcmplt <= '0';
                            ALUfunct <= "0000";
                            DRMUXSelt <= '0';
                            ACMUXSelt <= '0';
                            MemWRt <= '0';
                            MemREt <= '0';
                            RegBankaddrt <= IReg(9 downto 7); --changed
                            RegBankRWt <= '1'; --changed
                            RegBankImmValt <= "00000000";
                            RegBankImmEnt <= '0';
                            FGInRSTt <= '1';
                            FGOnRSTt <= '1';
                            nx_state <= T0;
                            when others =>
                        end case;
                    else -- immediate instruction
                        case (ImmInstOpcode) is
                            when "001" => -- ADDI
                                ArbiterSELt <= "000";
                                ARnRSTt <= '1';
                                PCnRSTt <= '1';
                                DRnRSTt <= '1';
                                EnRSTt <= '1';
                                ACnRSTt <= '1';
                                INPRnRSTt <= '1';
                                IRnRSTt <= '1';
                                RegBanknRSTt <= '1';
                                OUTRnRSTt <= '1';
                                ARLDt <= '0';
                                PCLDt <= '0';
                                DRLDt <= '0';
                                ACLDt <= '1'; --changed
                                INPRLDt <= '0';
                                IRLDt <= '0';
                                OUTRLDt <= '0';
                                ARInct <= '0';
                                PCInct <= '0';
                                DRInct <= '0';
                                ACInct <= '0';
                                INPRInct <= '0';
                                IRInct <= '0';
                                OUTRInct <= '0';
                                Ecmplt <= '0';
                                ACcmplt <= '0';
                                ALUfunct <= "0000"; --changed
                                DRMUXSelt <= '0'; --changed
                                ACMUXSelt <= '0'; --changed
                                MemWRt <= '0';
                                MemREt <= '0';
                                RegBankaddrt <= IReg(10 downto 8); --changed
                                RegBankRWt <= '0'; --changed
                                RegBankImmValt <= "00000000";
                                RegBankImmEnt <= '0';
                                FGInRSTt <= '1';
                                FGOnRSTt <= '1';
                                nx_state <= T6;
                            when others =>
                        end case;
                    end if;
                end if;
            when T6 =>
                ArbiterSELt <= "001"; --changed
                ARnRSTt <= '1';
                PCnRSTt <= '1';
                DRnRSTt <= '1';
                EnRSTt <= '1';
                ACnRSTt <= '1';
                INPRnRSTt <= '1';
                IRnRSTt <= '1';
                RegBanknRSTt <= '1';
                OUTRnRSTt <= '1';
                ARLDt <= '0';
                PCLDt <= '0';
                DRLDt <= '0';
                ACLDt <= '0';
                INPRLDt <= '0';
                IRLDt <= '0';
                OUTRLDt <= '0';
                ARInct <= '0';
                PCInct <= '0';
                DRInct <= '0';
                ACInct <= '0';
                INPRInct <= '0';
                IRInct <= '0';
                OUTRInct <= '0';
                Ecmplt <= '0';
                ACcmplt <= '0';
                ALUfunct <= "0000";
                DRMUXSelt <= '0';
                ACMUXSelt <= '0';
                MemWRt <= '0';
                MemREt <= '0';
                RegBankaddrt <= IReg(10 downto 8); --changed
                RegBankRWt <= '1'; --changed
                RegBankImmValt <= "00000000";
                RegBankImmEnt <= '0';
                FGInRSTt <= '1';
                FGOnRSTt <= '1';
                nx_state <= T6;
            when others =>
        end case;
    end process;

    process (pr_state, nRST, ArbiterSELt, ARnRSTt, PCnRSTt, DRnRSTt, EnRSTt, ACnRSTt, INPRnRSTt, IRnRSTt, RegBanknRSTt, OUTRnRSTt, ARLDt, PCLDt, DRLDt, ACLDt, INPRLDt, IRLDt, OUTRLDt, ARInct, PCInct, DRInct, ACInct, INPRInct, IRInct, OUTRInct, Ecmplt, ACcmplt, ALUfunct, DRMUXSelt, ACMUXSelt, MemWRt, MemREt, RegBankaddrt, RegBankRWt, RegBankImmValt, RegBankImmEnt, FGInRSTt, FGOnRSTt)
    begin
        if (nRST = '0') then
            ArbiterSEL <= "000";
            ARnRST <= '0';
            PCnRST <= '0';
            DRnRST <= '0';
            EnRST <= '0';
            ACnRST <= '0';
            INPRnRST <= '0';
            IRnRST <= '0';
            RegBanknRST <= '0';
            OUTRnRST <= '0';
            ARLD <= '0';
            PCLD <= '0';
            DRLD <= '0';
            ACLD <= '0';
            INPRLD <= '0';
            IRLD <= '0';
            OUTRLD <= '0';
            ARInc <= '0';
            PCInc <= '0';
            DRInc <= '0';
            ACInc <= '0';
            INPRInc <= '0';
            IRInc <= '0';
            OUTRInc <= '0';
            Ecmpl <= '0';
            ACcmpl <= '0';
            ALUfunc <= "0000";
            DRMUXSel <= '0';
            ACMUXSel <= '0';
            MemWR <= '0';
            MemRE <= '0';
            RegBankaddr <= "000";
            RegBankRW <= '0';
            RegBankImmVal <= "00000000";
            RegBankImmEn <= '0';
            FGInRST <= '1';
            FGOnRST <= '1';
            RInt <= '0';
        else
            ArbiterSEL <= ArbiterSELt;
            ARnRST <= ARnRSTt;
            PCnRST <= PCnRSTt;
            DRnRST <= DRnRSTt;
            EnRST <= EnRSTt;
            ACnRST <= ACnRSTt;
            INPRnRST <= INPRnRSTt;
            IRnRST <= IRnRSTt;
            RegBanknRST <= RegBanknRSTt;
            OUTRnRST <= OUTRnRSTt;
            ARLD <= ARLDt;
            PCLD <= PCLDt;
            DRLD <= DRLDt;
            ACLD <= ACLDt;
            INPRLD <= INPRLDt;
            IRLD <= IRLDt;
            OUTRLD <= OUTRLDt;
            ARInc <= ARInct;
            PCInc <= PCInct;
            DRInc <= DRInct;
            ACInc <= ACInct;
            INPRInc <= INPRInct;
            IRInc <= IRInct;
            OUTRInc <= OUTRInct;
            Ecmpl <= Ecmplt;
            ACcmpl <= ACcmplt;
            ALUfunc <= ALUfunct;
            DRMUXSel <= DRMUXSelt;
            ACMUXSel <= ACMUXSelt;
            MemWR <= MemWRt;
            MemRE <= MemREt;
            RegBankaddr <= RegBankaddrt;
            RegBankRW <= RegBankRWt;
            RegBankImmVal <= RegBankImmValt;
            RegBankImmEn <= RegBankImmEnt;
            FGInRST <= FGInRSTt;
            FGOnRST <= FGOnRSTt;
        end if;
    end process;

end Behavioral;

