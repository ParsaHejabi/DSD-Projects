-- $Id: prim.vhd,v 1.16 2001/10/16 18:40:26 pearl Exp pearl $
LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
LIBRARY IEEE;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;

package prim is

CONSTANT DefCombSpikeMsgOn : BOOLEAN := true;
CONSTANT DefCombSpikeXOn   : BOOLEAN := true;
CONSTANT DefSeqMsgOn       : BOOLEAN := true;
CONSTANT DefSeqXOn         : BOOLEAN := true;

CONSTANT DefDummyDelay      : VitalDelayType := 1.00 ns;
CONSTANT DefDummySetup      : VitalDelayType := 1.00 ns;
CONSTANT DefDummyHold       : VitalDelayType := 0.50 ns;
CONSTANT DefDummyWidth      : VitalDelayType := 1.00 ns;
CONSTANT DefDummyRecovery   : VitalDelayType := 1.00 ns;
CONSTANT DefDummyRecoverySR : VitalDelayType := 1.00 ns;
CONSTANT DefDummyRemoval    : VitalDelayType := 1.00 ns;
CONSTANT DefDummyIpd        : VitalDelayType := 0.00 ns;
CONSTANT DefDummyIsd        : VitalDelayType := 0.00 ns;
CONSTANT DefDummyIcd        : VitalDelayType := 0.00 ns;

CONSTANT udp_rfrd : VitalStateTableType (1 TO 5, 1 TO 4) := (
--      NOT,    IN      Q(t)   Q(t+1)
     (  'X',    '-',    '-',    'X'  ),
     (  '-',    '0',    '-',    '1'  ),
     (  '-',    '1',    '-',    '0'  ),
     (  '-',    '-',    '1',    '1'  ),
     (  '-',    '-',    '0',    '0'  ));

CONSTANT udp_dff : VitalStateTableType (1 TO 21, 1 TO 7) := (
--    NOTIFIER   D      CLK     RN       S      Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '0',    '-',    '1'  ),
     (  '-',    '-',    '-',    '0',    '1',    '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '1',    '-',    '0'  ),
     (  '-',    '1',    '/',    '1',    '-',    '-',    '1'  ),
     (  '-',    '1',    '*',    '1',    '-',    '1',    '1'  ),
     (  '-',    '0',    '*',    '-',    '1',    '0',    '0'  ),
     (  '-',    '-',    '\',    '-',    '-',    '-',    'S'  ),
     (  '-',    '*',    'B',    '-',    '-',    '-',    'S'  ),
     (  '-',    '-',    'B',    '1',    '*',    '1',    '1'  ),
     (  '-',    '1',    'X',    '1',    '*',    '1',    '1'  ),
     (  '-',    '-',    'B',    '*',    '1',    '0',    '0'  ),
     (  '-',    '0',    'X',    '*',    '1',    '0',    '0'  ),
     (  '-',    'B',    'r',    '-',    '-',    '-',    'X'  ),
     (  '-',    '/',    'X',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '*',    '-',    'X'  ),
     (  '-',    '-',    '-',    '*',    '-',    '-',    'X'  ),
     (  '-',    '-',    'f',    '-',    '-',    '-',    'X'  ),
     (  '-',    '\',    'X',    '1',    '-',    '-',    'X'  ),
     (  '-',    'B',    'X',    '-',    '-',    '-',    'S'  ),
     (  '-',    '-',    'S',    '-',    '-',    '-',    'S'  ));

CONSTANT udp_jkff : VitalStateTableType (1 TO 30, 1 TO 8) := (
--    NOTIFIER   J       K      CK       RN      SN     Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '-',    '0',    '-',    '1'  ),
     (  '-',    '-',    '-',    '-',    '0',    '1',    '-',    '0'  ),
     (  '-',    '0',    '0',    '/',    '1',    '1',    '-',    'S'  ),  
     (  '-',    '0',    '1',    '/',    '-',    '1',    '-',    '0'  ), 
     (  '-',    '1',    '0',    '/',    '1',    '-',    '-',    '1'  ),
     (  '-',    '-',    '1',    '/',    '-',    '1',    '1',    '0'  ),
     (  '-',    '1',    '-',    '/',    '1',    '-',    '0',    '1'  ),
     (  '-',    '-',    '0',    '*',    '1',    '-',    '1',    '1'  ),
     (  '-',    '0',    '-',    '*',    '-',    '1',    '0',    '0'  ),
     (  '-',    '-',    '-',    '\',    '-',    '-',    '-',    'S'  ),
     (  '-',    '*',    '-',    'B',    '-',    '-',    '-',    'S'  ),
     (  '-',    '*',    '0',    '-',    '1',    '-',    '1',    '1'  ),
     (  '-',    '-',    '*',    'B',    '-',    '-',    '-',    'S'  ),
     (  '-',    '0',    '*',    '-',    '-',    '1',    '0',    '0'  ),
     (  '-',    '-',    '-',    'B',    '1',    '*',    '1',    '1'  ),
     (  '-',    '-',    '0',    'X',    '1',    '*',    '1',    '1'  ),
     (  '-',    '-',    '-',    'B',    '*',    '1',    '0',    '0'  ),
     (  '-',    '0',    '-',    'X',    '*',    '1',    '0',    '0'  ),
     (  '-',    '0',    'S',    '-',    '-',    '1',    '0',    '0'  ),
     (  '-',    '0',    'X',    '-',    'X',    '1',    '0',    '0'  ),
     (  '-',    'S',    '0',    '-',    '1',    '-',    '1',    '1'  ),
     (  '-',    'X',    '0',    '-',    '1',    'X',    '1',    '1'  ),
     (  '-',    '-',    '-',    '-',    '-',    '*',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '*',    '-',    '-',    'X'  ),
     (  '-',    '*',    '-',    'X',    '1',    '1',    '-',    'X'  ),
     (  '-',    '-',    '*',    'X',    '1',    '1',    '-',    'X'  ),
     (  '-',    '-',    '-',    '*',    '1',    '1',    '-',    'X'  ),
     (  '-',    '-',    '-',    'X',    '1',    '1',    '-',    'S'  ),
     (  '-',    '-',    '-',    'S',    '-',    '-',    '-',    'S'  ));

CONSTANT udp_sjkff : VitalStateTableType (1 TO 42, 1 TO 10) := (
--    NOTIFIER   SE    SI    J      K     CK      RN     SN    Q(t)   Q(t+1)
     (  'X',    '-',  '-',  '-',   '-',   '-',   '-',   '-',   '-',    'X'  ),
     (  '-',    '-',  '-',  '-',   '-',   '-',   '-',   '0',   '-',    '1'  ),
     (  '-',    '-',  '-',  '-',   '-',   '-',   '0',   '1',   '-',    '0'  ),
     (  '-',    '0',  '-',  '0',   '0',   '/',   '1',   '1',   '-',    'S'  ),  
     (  '-',    '0',  '-',  '0',   '1',   '/',   '-',   '1',   '-',    '0'  ), 
     (  '-',    '0',  '-',  '1',   '0',   '/',   '1',   '-',   '-',    '1'  ), 
     (  '-',    '0',  '-',  '1',   '1',   '/',   '1',   '1',   '1',    '0'  ), 
     (  '-',    '0',  '-',  '1',   '1',   '/',   '1',   '1',   '0',    '1'  ),
     (  '-',    '1',  '0',  '-',   '-',   '/',   '-',   '1',   '-',    '0'  ),
     (  '-',    '1',  '1',  '-',   '-',   '/',   '1',   '-',   '-',    '1'  ),
     (  '-',    '-',  '1',  '1',   '0',   '/',   '1',   '-',   '-',    '1'  ),
     (  '-',    '-',  '0',  '0',   '1',   '/',   '-',   '1',   '-',    '0'  ),
     (  '-',    '0',  '-',  '-',   '0',   '-',   '1',   '-',   '1',    '1'  ),
     (  '-',    '1',  '1',  '-',   '-',   '-',   '1',   '-',   '1',    '1'  ),
     (  '-',    '0',  '-',  '0',   '-',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '0',  '-',  '0',   '0',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '0',  '-',  '0',   '0',   '-',   '1',   '-',   '1',    '1'  ),
     (  '-',    '0',  '-',  '0',   '0',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '0',  '-',  '0',   '-',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '1',  '0',  '-',   '-',   '-',   '-',   '1',   '0',    'S'  ),
     (  '-',    '-',  '-',  '-',   '-',   '\',   '-',   '-',   '-',    'S'  ),
     (  '-',    '*',  '-',  '-',   '-',   'B',   '-',   '-',   '-',    'S'  ),
     (  '-',    '-',  '*',  '-',   '-',   'B',   '-',   '-',   '-',    'S'  ),
     (  '-',    '-',  '-',  '*',   '-',   'B',   '-',   '-',   '-',    'S'  ),
     (  '-',    '-',  '1',  '-',   '0',   '-',   '1',   '-',   '1',    '1'  ),
     (  '-',    '-',  '0',  '0',   '-',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '0',  '-',  '*',   '0',   '-',   '1',   '-',   '1',    '1'  ),
     (  '-',    '-',  '-',  '-',   '*',   'B',   '-',   '-',   '-',    'S'  ),
     (  '-',    '0',  '-',  '0',   '*',   '-',   '-',   '1',   '0',    '0'  ),
     (  '-',    '0',  '*',  '-',   '-',   '-',   '-',   '-',   '-',    'S'  ),
     (  '-',    '1',  '-',  '*',   '-',   '-',   '-',   '-',   '-',    'S'  ),
     (  '-',    '1',  '-',  '-',   '*',   '-',   '-',   '-',   '-',    'S'  ),
     (  '-',    '-',  '-',  '-',   '-',   'B',   '0',   'X',   '-',    'X'  ),
     (  '-',    '-',  '-',  '-',   '-',   'B',   'X',   'X',   '-',    'X'  ),
     (  '-',    '-',  '-',  '-',   '-',   'B',   'X',   '1',   '1',    'X'  ),
     (  '-',    '-',  '-',  '-',   '-',   'B',   '1',   'X',   '0',    'X'  ),
     (  '-',    '0',  '-',  '-',   '0',   '-',   '1',   '*',   '1',    'S'  ),
     (  '-',    '1',  '1',  '-',   '-',   '-',   '1',   '*',   '1',    'S'  ),
     (  '-',    '-',  '-',  '-',   '-',   'B',   '*',   '1',   '0',    'S'  ),
     (  '-',    '0',  '-',  '0',   '-',   '-',   '*',   '1',   '0',    'S'  ),
     (  '-',    '1',  '0',  '-',   '-',   '-',   '*',   '1',   '0',    'S'  ),
     (  '-',    '-',  '-',  '-',   '-',   'S',   '-',   '-',    '-',   'S'  ));


CONSTANT udp_xgen4 : VitalTruthTableType (1 TO 12, 1 TO 10) := (
     (  '1',    '1',    '-',  '-',  '-',  '-',  '-',  '-',  '-',    'X'  ),
     (  '0',    '0',    '-',  '-',  '-',  '-',  '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '1',  '1',  '-',  '-',  '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '0',  '0',  '-',  '-',  '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '-',  '-',  '1',  '1',  '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '-',  '-',  '0',  '0',  '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '-',  '-',  '-',  '-',  '1',  '1',  '-',    'X'  ),
     (  '-',    '-',    '-',  '-',  '-',  '-',  '0',  '0',  '-',    'X'  ),
     (  '0',    '1',    '-',  '-',  '-',  '-',  '-',  '-',  '1',    '1'  ),
     (  '0',    '1',    '-',  '-',  '-',  '-',  '-',  '-',  '0',    '0'  ),
     (  '1',    '0',    '-',  '-',  '-',  '-',  '-',  '-',  '1',    '1'  ),
     (  '1',    '0',    '-',  '-',  '-',  '-',  '-',  '-',  '0',    '0'  ));

CONSTANT udp_xgen : VitalTruthTableType (1 TO 6, 1 TO 4) := (
     (  '1',    '1',    '-',    'X'  ),
     (  '0',    '0',    '-',    'X'  ),
     (  '0',    '1',    '1',    '1'  ),
     (  '0',    '1',    '0',    '0'  ),
     (  '1',    '0',    '1',    '1'  ),
     (  '1',    '0',    '0',    '0'  ));

CONSTANT udp_outrf : VitalTruthTableType (1 TO 5, 1 TO 4) := (
     (  '1',    '-',    '0',    '1'  ),
     (  '0',    '1',    '-',    '1'  ),
     (  '-',    '0',    '1',    '0'  ),
     (  '0',    '0',    '-',    '0'  ),
     (  '1',    '-',    '1',    '0'  ));

CONSTANT udp_mux : VitalTruthTableType (1 TO 6, 1 TO 4) := (
     (  '1',    '-',    '0',    '1'  ),
     (  '0',    '-',    '0',    '0'  ),
     (  '-',    '1',    '1',    '1'  ),
     (  '-',    '0',    '1',    '0'  ),
     (  '0',    '0',    'X',    '0'  ),
     (  '1',    '1',    'X',    '1'  )  );


CONSTANT udp_mux2 : VitalTruthTableType (1 TO 6, 1 TO 4) := (
     (  '1',    '-',    '0',    '1'  ),
     (  '0',    '-',    '0',    '0'  ),
     (  '-',    '1',    '1',    '1'  ),
     (  '-',    '0',    '1',    '0'  ),
     (  '0',    '0',    'X',    '0'  ),
     (  '1',    '1',    'X',    '1'  )  );


CONSTANT udp_mux4 : VitalTruthTableType (1 TO 18, 1 TO 7) := (
     (  '0',    '-',    '-',    '-',    '0',    '0',    '0'  ),
     (  '1',    '-',    '-',    '-',    '0',    '0',    '1'  ),
     (  '-',    '0',    '-',    '-',    '1',    '0',    '0'  ),
     (  '-',    '1',    '-',    '-',    '1',    '0',    '1'  ),
     (  '-',    '-',    '0',    '-',    '0',    '1',    '0'  ),
     (  '-',    '-',    '1',    '-',    '0',    '1',    '1'  ),
     (  '-',    '-',    '-',    '0',    '1',    '1',    '0'  ),
     (  '-',    '-',    '-',    '1',    '1',    '1',    '1'  ),
     (  '0',    '0',    '-',    '-',    'X',    '0',    '0'  ),
     (  '1',    '1',    '-',    '-',    'X',    '0',    '1'  ),
     (  '-',    '-',    '0',    '0',    'X',    '1',    '0'  ),
     (  '-',    '-',    '1',    '1',    'X',    '1',    '1'  ),
     (  '0',    '-',    '0',    '-',    '0',    'X',    '0'  ),
     (  '1',    '-',    '1',    '-',    '0',    'X',    '1'  ),
     (  '-',    '0',    '-',    '0',    '1',    'X',    '0'  ),
     (  '-',    '1',    '-',    '1',    '1',    'X',    '1'  ),
     (  '1',    '1',    '1',    '1',    'X',    'X',    '1'  ),
     (  '0',    '0',    '0',    '0',    'X',    'X',    '0'  )  );

CONSTANT udp_bmux : VitalTruthTableType (1 TO 14, 1 TO 6) := (
     (  '0',   '-',   '0',   '1',   '-',    '0' ),
     (  '1',   '-',   '0',   '-',   '0',    '1' ),
     (  '-',   '0',   '1',   '1',   '-',    '0' ),
     (  '-',   '1',   '1',   '-',   '0',    '1' ),
     (  '0',   '0',   '-',   '1',   '-',    '0' ),
     (  '1',   '1',   '-',   '-',   '0',    '1' ),
     (  '0',   '-',   '0',   '0',   '-',    '1' ),
     (  '1',   '-',   '0',   '-',   '1',    '0' ),
     (  '-',   '0',   '1',   '0',   '-',    '1' ),
     (  '-',   '1',   '1',   '-',   '1',    '0' ),
     (  '0',   '0',   '-',   '0',   '-',    '1' ),
     (  '1',   '1',   '-',   '-',   '1',    '0' ),
     (  '-',   '-',   '-',   '0',   '0',    '1' ),
     (  '-',   '-',   '-',   '1',   '1',    '0' ));

CONSTANT udp_bmx : VitalTruthTableType (1 TO 12, 1 TO 6) := (
     (  '0',   '1',   '1',   '-',   '-',    '0' ),
     (  '0',   '1',   '0',   '0',   '-',    '1' ),
     (  '0',   '1',   '0',   '1',   '-',    '0' ),
     (  '0',   '0',   '1',   '0',   '-',    '0' ),
     (  '0',   '0',   '1',   '1',   '-',    '1' ),
     (  '0',   '0',   '0',   '-',   '-',    '1' ),
     (  '1',   '1',   '1',   '-',   '-',    '0' ),
     (  '1',   '1',   '0',   '-',   '0',    '1' ),
     (  '1',   '1',   '0',   '-',   '1',    '0' ),
     (  '1',   '0',   '1',   '-',   '0',    '0' ),
     (  '1',   '0',   '1',   '-',   '1',    '1' ),
     (  '1',   '0',   '0',   '-',   '-',    '1' ));

CONSTANT udp_rslat_out : VitalStateTableType (1 TO 22, 1 TO 5) := (
     (  'X',    '-',    '-',    '-',    'X'  ),
     (  '-',    '\',    '0',    '-',    'S'  ),
     (  '-',    'v',    '0',    '-',    'S'  ),
     (  '-',    '0',    '\',    '-',    'S'  ),
     (  '-',    '0',    'v',    '-',    'S'  ),
     (  '-',    '/',    '0',    '-',    '0'  ),
     (  '-',    '^',    '0',    '-',    '0'  ),
     (  '-',    '1',    '-',    '-',    '0'  ),
     (  '-',    '\',    '1',    '-',    '1'  ),
     (  '-',    'v',    '1',    '-',    '1'  ),
     (  '-',    '0',    '/',    '-',    '1'  ),
     (  '-',    '0',    '^',    '-',    '1'  ),
     (  '-',    '/',    '1',    '-',    '0'  ),
     (  '-',    '^',    '1',    '-',    '0'  ),
     (  '-',    '\',    'X',    '1',    '1'  ),
     (  '-',    'v',    'X',    '1',    '1'  ),
     (  '-',    '0',    'r',    '1',    '1'  ),
     (  '-',    '0',    'f',    '1',    '1'  ),
     (  '-',    'r',    '0',    '0',    '0'  ),
     (  '-',    'f',    '0',    '0',    '0'  ),
     (  '-',    'X',    '\',    '0',    '0'  ),
     (  '-',    'X',    'v',    '0',    '0'  )  );


CONSTANT udp_rslat_out_n : VitalStateTableType (1 TO 22, 1 TO 5) := (
     (  'X',    '-',    '-',    '-',    'X'  ),
     (  '-',    '\',    '0',    '-',    'S'  ),
     (  '-',    'v',    '0',    '-',    'S'  ),
     (  '-',    '0',    '\',    '-',    'S'  ),
     (  '-',    '0',    'v',    '-',    'S'  ),
     (  '-',    '/',    '0',    '-',    '1'  ),
     (  '-',    '^',    '0',    '-',    '1'  ),
     (  '-',    '1',    '\',    '-',    '1'  ),
     (  '-',    '1',    'v',    '-',    '1'  ),
     (  '-',    '-',    '1',    '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '0'  ),
     (  '-',    '0',    '^',    '-',    '0'  ),
     (  '-',    '1',    '/',    '-',    '0'  ),
     (  '-',    '1',    '^',    '-',    '0'  ),
     (  '-',    '\',    'X',    '0',    '0'  ),
     (  '-',    'v',    'X',    '0',    '0'  ),
     (  '-',    '0',    'r',    '0',    '0'  ),
     (  '-',    '0',    'f',    '0',    '0'  ),
     (  '-',    'r',    '0',    '1',    '1'  ),
     (  '-',    'f',    '0',    '1',    '1'  ),
     (  '-',    'X',    '\',    '1',    '1'  ),
     (  '-',    'X',    'v',    '1',    '1'  )  );


CONSTANT udp_rslatn_out : VitalStateTableType (1 TO 22, 1 TO 5) := (
     (  'X',    '-',    '-',    '-',    'X'  ),
     (  '-',    '/',    '1',    '-',    'S'  ),
     (  '-',    '^',    '1',    '-',    'S'  ),
     (  '-',    '1',    '/',    '-',    'S'  ),
     (  '-',    '1',    '^',    '-',    'S'  ),
     (  '-',    '\',    '1',    '-',    '0'  ),
     (  '-',    'v',    '1',    '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '0'  ),
     (  '-',    '0',    '^',    '-',    '0'  ),
     (  '-',    '0',    '\',    '-',    '1'  ),
     (  '-',    '0',    'v',    '-',    '1'  ),
     (  '-',    '-',    '0',    '-',    '1'  ),
     (  '-',    '1',    '\',    '-',    '1'  ),
     (  '-',    '1',    'v',    '-',    '1'  ),
     (  '-',    '/',    'X',    '1',    '1'  ),
     (  '-',    '^',    'X',    '1',    '1'  ),
     (  '-',    '1',    'r',    '1',    '1'  ),
     (  '-',    '1',    'f',    '1',    '1'  ),
     (  '-',    'r',    '1',    '0',    '0'  ),
     (  '-',    'f',    '1',    '0',    '0'  ),
     (  '-',    'X',    '/',    '0',    '0'  ),
     (  '-',    'X',    '^',    '0',    '0'  )  );


CONSTANT udp_rslatn_out_n : VitalStateTableType (1 TO 22, 1 TO 5) := (
     (  'X',    '-',    '-',    '-',    'X'  ),
     (  '-',    '/',    '1',    '-',    'S'  ),
     (  '-',    '^',    '1',    '-',    'S'  ),
     (  '-',    '1',    '/',    '-',    'S'  ),
     (  '-',    '1',    '^',    '-',    'S'  ),
     (  '-',    '\',    '1',    '-',    '1'  ),
     (  '-',    'v',    '1',    '-',    '1'  ),
     (  '-',    '0',    '-',    '-',    '1'  ),
     (  '-',    '/',    '0',    '-',    '0'  ),
     (  '-',    '^',    '0',    '-',    '0'  ),
     (  '-',    '\',    '0',    '-',    '1'  ),
     (  '-',    'v',    '0',    '-',    '1'  ),
     (  '-',    '1',    '\',    '-',    '0'  ),
     (  '-',    '1',    'v',    '-',    '0'  ),
     (  '-',    '/',    'X',    '0',    '0'  ),
     (  '-',    '^',    'X',    '0',    '0'  ),
     (  '-',    '1',    'r',    '0',    '0'  ),
     (  '-',    '1',    'f',    '0',    '0'  ),
     (  '-',    'r',    '1',    '1',    '1'  ),
     (  '-',    'f',    '1',    '1',    '1'  ),
     (  '-',    'X',    '/',    '1',    '1'  ),
     (  '-',    'X',    '^',    '1',    '1'  )  );

CONSTANT udp_tlatrf : VitalStateTableType (1 TO 6, 1 TO 6) := (
--      NOT      D       G      GN       Q(t)  Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '1',    '1',    '0',    '-',    '0'  ), 
     (  '-',    '0',    '1',    '0',    '-',    '1'  ), 
     (  '-',    '0',    '-',    '-',    '1',    '1'  ), 
     (  '-',    '1',    '-',    '-',    '0',    '0'  ), 
     (  '-',    '-',    '0',    '1',    '-',    'S'  ));

CONSTANT udp_tlatrf2 : VitalStateTableType (1 TO 12, 1 TO 7) := (
--      NOT      D1      G1      D2      G2      Q(t)  Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',     '-',  'X'  ),
     (  '-',    '1',    '1',    '-',    '0',     '-',  '1'  ), 
     (  '-',    '0',    '1',    '-',    '0',     '-',  '0'  ), 
     (  '-',    '-',    '0',    '0',    '1',     '-',  '0'  ), 
     (  '-',    '-',    '0',    '1',    '1',     '-',  '1'  ), 
     (  '-',    '1',    '1',    '1',    '1',     '-',  '1'  ), 
     (  '-',    '0',    '1',    '0',    '1',     '-',  '0'  ), 
     (  '-',    '0',    'X',    '-',    '0',     '0',  '0'  ), 
     (  '-',    '1',    'X',    '-',    '0',     '1',  '1'  ), 
     (  '-',    '-',    '0',    '0',    'X',     '0',  '0'  ), 
     (  '-',    '-',    '0',    '1',    'X',     '1',  '1'  ), 
     (  '-',    '-',    '0',    '-',    '0',     '-',  'S'  ));


CONSTANT udp_tlat : VitalStateTableType (1 TO 20, 1 TO 7) := (
--      NOT      D       G       R       S      Q(t)  Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '0',    '-',    '1'  ),
     (  '-',    '-',    '-',    '0',    '1',    '-',    '0'  ),
     (  '-',    '1',    '0',    '1',    '-',    '-',    '1'  ), 
     (  '-',    '0',    '0',    '-',    '1',    '-',    '0'  ), 
     (  '-',    '1',    '*',    '1',    '-',    '1',    '1'  ),
     (  '-',    '0',    '*',    '-',    '1',    '0',    '0'  ),
     (  '-',    '*',    '1',    '-',    '-',    '-',    'S'  ),
     (  '-',    '-',    '1',    '1',    '*',    '1',    '1'  ),
     (  '-',    '1',    '-',    '1',    '*',    '1',    '1'  ),
     (  '-',    '-',    '1',    '*',    '1',    '0',    '0'  ),
     (  '-',    '0',    '-',    '*',    '1',    '0',    '0'  ),
     (  '-',    '0',    '-',    '-',    '1',    '0',    '0'  ),
     (  '-',    '1',    '-',    '1',    '-',    '1',    '1'  ),
     (  '-',    '*',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '*',    '-',    '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '*',    '-',    'X'  ),
     (  '-',    'B',    'f',    '1',    '1',    '-',    'X'  ),
     (  '-',    'B',    'X',    '1',    '1',    '-',    'S'  ),
     (  '-',    '-',    'S',    '-',    '-',    '-',    'S'  ) ); 

CONSTANT udp_etlat : VitalStateTableType (1 TO 31, 1 TO 8) := (
--      NOT      D       G       R       S     E    Q(t)  Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',  '-',  '-',    'X'  ),
     (  '-',    '1',    '0',    '1',    '1',  '1',  '-',    '1'  ),
     (  '-',    '0',    '0',    '1',    '1',  '1',  '-',    '0'  ),
     (  '-',    '-',    '/',    '1',    '1',  '0',  '-',    'S'  ),
     (  '-',    '-',    '1',    '1',    '1',  '\',  '-',    'S'  ),
     (  '-',    '-',    '\',    '1',    '1',  '0',  '-',    'S'  ),
     (  '-',    '-',    '1',    '1',    '1',  '/',  '-',    'S'  ),
     (  '-',    '0',    '/',    '1',    '1',  '1',  '-',    '0'  ),
     (  '-',    '1',    '/',    '1',    '1',  '1',  '-',    '1'  ),
     (  '-',    '0',    '0',    '1',    '1',  '\',  '-',    '0'  ),
     (  '-',    '1',    '0',    '1',    '1',  '\',  '-',    '1'  ),
     (  '-',    '1',    '*',    '1',    '-',  '1',  '1',    '1'  ),
     (  '-',    '0',    '*',    '-',    '1',  '1',  '0',    '0'  ),
     (  '-',    '1',    '0',    '1',    '-',  '*',  '1',    '1'  ),
     (  '-',    '0',    '0',    '-',    '1',  '*',  '0',    '0'  ),
     (  '-',    '*',    '1',    '-',    '-',  '-',  '-',    'S'  ),
     (  '-',    '*',    '-',    '-',    '-',  '0',  '-',    'S'  ),
     (  '-',    '-',    '-',    '-',    '0',  '-',  '-',    '1'  ),
     (  '-',    '-',    '1',    '1',    '*',  '-',  '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '*',  '0',  '1',    '1'  ),
     (  '-',    '1',    '-',    '1',    '*',  '-',  '1',    '1'  ),
     (  '-',    '-',    '-',    '0',    '1',  '-',  '-',    '0'  ),
     (  '-',    '-',    '1',    '*',    '1',  '-',  '0',    '0'  ),
     (  '-',    '-',    '-',    '*',    '1',  '0',  '0',    '0'  ),
     (  '-',    '0',    '-',    '*',    '1',  '-',  '0',    '0'  ),
 
     --(  '-',    '0',    '-',    '-',    '1',  '1',  '0',    '0'  ),
     --(  '-',    '1',    '-',    '1',    '-',  '1',  '1',    '1'  ),
     (  '-',    '*',    '-',    '-',    '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '-',    '*',    '-',  '-',  '-',    'X'  ),
     (  '-',    '-',    '-',    '-',    '*',  '-',  '-',    'X'  ),
     (  '-',    'B',    'f',    '1',    '1',  '-',  '-',    'X'  ),
     (  '-',    'B',    'X',    '1',    '1',  '-',  '-',    'S'  ),
     (  '-',    '-',    'S',    '-',    '-',  '-',  '-',    'S'  ) ); 


CONSTANT udp_edfft : VitalStateTableType (1 TO 23, 1 TO 8) := (
--    NOTIFIER   D      CLK     RN       S      EN    Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',    '-',    'X'  ),
     (  '-',    '-',    '/',    '0',    '1',    '-',    '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '1',    '1',    '-',    '0'  ),
     (  '-',    '-',    '/',    '-',    '0',    '-',    '-',    '1'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',    '-',    '1'  ),
     (  '-',    '-',    '-',    '1',    '1',    '0',    '-',    'S'  ),
     (  '-',    '1',    '*',    '1',    '-',    '-',    '1',    '1'  ),
     (  '-',    '-',    '*',    '-',    '0',    '-',    '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '-',    '0',    '1',    '1'  ),
     (  '-',    '0',    '*',    '-',    '1',    '-',    '0',    '0'  ),
     (  '-',    '-',    '*',    '0',    '1',    '-',    '0',    '0'  ),
     (  '-',    '-',    '-',    '-',    '1',    '0',    '0',    '0'  ),
     (  '-',    '-',    '\',    '-',    '-',    '-',    '-',    'S'  ),
     (  '-',    '-',    'v',    '-',    '-',    '-',    '-',    'S'  ),
     (  '-',    '*',    'B',    '-',    '-',    '-',    '-',    'S'  ),
     (  '-',    '1',    'X',    '1',    '-',    '-',    '1',    '1'  ),
     (  '-',    '0',    'X',    '-',    '1',    '-',    '0',    '0'  ),
     (  '-',    '-',    'B',    '-',    '-',    '*',    '-',    'S'  ),
     (  '-',    '-',    'B',    '*',    '-',    '-',    '-',    'S'  ),
     (  '-',    '-',    'X',    '0',    '1',    '-',    '0',    '0'  ),
     (  '-',    '-',    'B',    '-',    '*',    '-',    '-',    'S'  ),
     (  '-',    '-',    'X',    '-',    '0',    '-',    '1',    '1'  ),
     (  '-',    '-',    'S',    '-',    '-',    '-',    '-',    'S'  ));

CONSTANT udp_sedfft : VitalStateTableType (1 TO 53, 1 TO 10) := (
--    NOTIFIER   D      CLK     RN       S      EN    SI   SE   Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',  '-', '-', '-',    'X'  ),
     (  '-',    '-',    '/',    '-',    '-',    '-',  '0', '1', '-',    '0'  ),
     (  '-',    '-',    '/',    '-',    '-',    '-',  '1', '1', '-',    '1'  ),
     (  '-',    '-',    'B',    '-',    '-',    '-',  '-', '*', '-',    'S'  ),
     (  '-',    '-',    'B',    '-',    '-',    '-',  '*', '-', '-',    'S'  ),
     (  '-',    '-',    '\',    '-',    '-',    '-',  '-', '-',  '-',   'S'  ),
     (  '-',    '-',    'v',    '-',    '-',    '-',  '-', '-',  '-',   'S'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',  '1', '-', '-',    '1'  ),
     (  '-',    '0',    '/',    '-',    '1',    '1',  '0', '-', '-',    '0'  ),
     (  '-',    '1',    '/',    '1',    '-',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '0',    '/',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '-',    '/',    '-',    '0',    '-',  '1', '-', '-',    '1'  ),
     (  '-',    '-',    '/',    '0',    '1',    '-',  '0', '-', '-',    '0'  ),
     (  '-',    '-',    'X',    '-',    '-',    '-',  '0', '1', '0',    'S'  ),
     (  '-',    '-',    'X',    '-',    '-',    '-',  '1', '1', '1',    'S'  ),
     (  '-',    '-',    'X',    '-',    '0',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    'X',    '0',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '1',    'X',    '1',    '-',    '1',  '1', '-', '1',    '1'  ),
     (  '-',    '0',    'X',    '-',    '1',    '1',  '0', '-', '0',    '0'  ),
     (  '-',    '-',    '-',    '-',    '1',    '0',  '-', '0', '0',    '0'  ), -- new
     (  '-',    '-',    '-',    '-',    '1',    '0',  '0', '-', '0',    '0'  ), -- new
     (  '-',    '-',    '-',    '1',    '1',    '0',  '1', '-', '1',    '1'  ), -- new
     (  '-',    '-',    '-',    '-',    '1',    '0',  '-', '0', '0',    '0'  ), -- new
     (  '-',    '-',    '-',    '1',    '-',    '0',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '1',    '0',  '-', '0', '-',    'S'  ), -- new
     (  '-',    '-',    '/',    '0',    '1',    '-',  '-', '0', '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '1',    '1',  '-', '0', '-',    '0'  ),
     (  '-',    '-',    '/',    '-',    '0',    '-',  '-', '0', '-',    '1'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',  '-', '0', '-',    '1'  ),
     (  '-',    '-',    '/',    '1',    '1',    '0',  '-', '0', '-',    'S'  ),
     (  '-',    '-',    '-',    '-',    '-',    '-',  '0', '1', '0',    '0'  ),
     (  '-',    '-',    '-',    '0',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '0',    '-',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '1',    '-',    '1',    '-',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '0',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '-',    '-',    '-',    '-',  '1', '1', '1',    '1'  ),
     (  '-',    '1',    '*',    '1',    '-',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '*',    '-',    '0',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '*',    '-',    '0',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '1',    '*',    '1',    '-',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '*',    '0',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    '*',    '0',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '0',    '*',    '-',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '0',    '*',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '*',    'B',    '-',    '-',    '-',  '-', '-', '-',    'S'  ),
     (  '-',    '1',    'X',    '1',    '-',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '0',    'X',    '-',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    'B',    '-',    '-',    '*',  '-', '-', '-',    'S'  ),
     (  '-',    '-',    'B',    '*',    '-',    '-',  '-', '-', '-',    'S'  ),
     (  '-',    '-',    'X',    '0',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    'B',    '-',    '*',    '-',  '-', '-', '-',    'S'  ),
     (  '-',    '-',    'X',    '-',    '0',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    'S',    '-',    '-',    '-',  '-', '-', '-',    'S'  ));

CONSTANT udp_edff : VitalStateTableType (1 TO 21, 1 TO 8) := (
--    NOTIFIER   D      CLK     RN       S      EN    Q(t)   Q(t+1)
       (  'X',    '-',    '-',    '-',    '-',    '-',    '-',    'X'  ),
       (  '-',    '-',    '-',    '-',    '0',    '-',    '-',    '1'  ),
       (  '-',    '-',    '-',    '0',    '1',    '-',    '-',    '0'  ),
       (  '-',    '0',    '/',    '-',    '1',    '1',    '-',    '0'  ),
       (  '-',    '1',    '/',    '1',    '-',    '1',    '-',    '1'  ),
       (  '-',    '-',    '*',    '-',    '-',    '0',    '-',    'S'  ),
       (  '-',    '1',    '*',    '1',    '-',    '-',    '1',    '1'  ),
       (  '-',    '0',    '*',    '-',    '1',    '-',    '0',    '0'  ),
       (  '-',    '-',    '\',    '-',    '-',    '-',    '-',    'S'  ),
       (  '-',    '*',    'B',    '-',    '-',    '-',    '-',    'S'  ),
       (  '-',    '1',    'X',    '1',    '-',    '-',    '1',    '1'  ),
       (  '-',    '0',    'X',    '-',    '1',    '-',    '0',    '0'  ),
       (  '-',    '-',    'B',    '-',    '-',    '*',    '-',    'S'  ),
       (  '-',    '-',    'X',    '1',    '1',    '0',    '-',    'S'  ),
       (  '-',    '-',    'X',    'X',    '1',    '0',    '0',    '0'  ),
       (  '-',    '-',    'X',    '1',    'X',    '0',    '1',    '1'  ),
       (  '-',    '-',    'B',    '1',    '*',    '-',    '1',    '1'  ),
       (  '-',    '-',    'B',    '*',    '1',    '-',    '0',    '0'  ),
       (  '-',    '-',    '-',    '-',    '*',    '-',    '-',    'X'  ),
       (  '-',    '-',    '-',    '*',    '-',    '-',    '-',    'X'  ),
       (  '-',    '-',    'S',    '-',    '-',    '-',    '-',    'S'  ));

CONSTANT udp_sedff : VitalStateTableType (1 TO 42, 1 TO 10) := ( 
--    NOTIFIER   D      CLK     RN       S      EN    SI   SE   Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',  '-', '-', '-',    'X'  ),
     (  '-',    '-',    '-',    '0',    '1',    '-',  '-', '-', '-',    '0'  ),
     (  '-',    '-',    '/',    '-',    '-',    '-',  '0', '1', '-',    '0'  ),
     (  '-',    '-',    '/',    '1',    '-',    '-',  '1', '1', '-',    '1'  ),
     (  '-',    '-',    'B',    '*',    '1',    '-',  '-', '-', '0',    '0'  ),
     (  '-',    '-',    'B',    'p',    '1',    '-',  '-', '-', '1',    'X'  ),
     (  '-',    '-',    'B',    'n',    '1',    '-',  '-', '-', '1',    'X'  ),
     (  '-',    '*',    'B',    '-',    '-',    '-',  '-', '-', '-',    'S'  ),
     (  '-',    '*',    '-',    '-',    '-',    '0',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    'B',    '1',    '*',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    'B',    '-',    '-',    '*',  '-', '-', '-',    'S'  ),
     (  '-',    '-',    'B',    '-',    '-',    '-',  '-', '*', '-',    'S'  ),
     (  '-',    '-',    'B',    '-',    '-',    '-',  '*', '-', '-',    'S'  ),
     (  '-',    '-',    '\',    '-',    '-',    '-',  '-', '-',  '-',   'S'  ),
     (  '-',    '-',    '-',    '1',    '-',    '0',  '-', '0',  '1',   '1'  ),
     (  '-',    '-',    '-',    '-',    '1',    '0',  '-', '0',  '0',   '0'  ),
     (  '-',    '-',    'X',    '-',    '-',    '-',  '0', '1', '0',    '0'  ),
     (  '-',    '1',    '-',    '1',    '-',    '-',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '-',    '-',  '1', '1', '1',    '1'  ),
     (  '-',    '0',    '-',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),
     (  '-',    '-',    '-',    '-',    '1',    '-',  '0', '1', '0',    '0'  ),
     (  '-',    '-',    'X',    '1',    '-',    '-',  '1', '1', '1',    '1'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',  '1', '-', '-',    '1'  ),
     (  '-',    '0',    '/',    '-',    '1',    '1',  '0', '-', '-',    '0'  ),
     (  '-',    '1',    'X',    '1',    '-',    '1',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    'X',    '1',    '-',    '0',  '1', '-', '1',    '1'  ),
     (  '-',    '0',    'X',    '-',    '1',    '1',  '0', '-', '0',    '0'  ),
     (  '-',    '-',    'X',    '-',    '1',    '0',  '0', '-', '0',    '0'  ),
     (  '-',    '0',    '/',    '-',    '1',    '1',  '-', '0', '-',    '0'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',  '-', '0', '-',    '1'  ),
     (  '-',    '-',    '*',    '-',    '1',    '0',  '0', '-', '0',    '0'  ),
     (  '-',    '-',    '*',    '-',    '1',    '0',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    '*',    '1',    '-',    '0',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '/',    '-',    '-',    '0',  '-', '0', '-',    'S'  ),
     (  '-',    '1',    '*',    '1',    '-',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '*',    '1',    '-',    '0',  '-', '0', '1',    '1'  ),
     (  '-',    '0',    '*',    '-',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '1',    'X',    '1',    '-',    '-',  '-', '0', '1',    '1'  ),
     (  '-',    '0',    'X',    '-',    '1',    '-',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    'X',    '1',    '1',    '0',  '-', '0', '-',    'S'  ),
     (  '-',    '-',    '-',    '1',    '0',    '-',  '-', '-', '-',    '1'  ),
     (  '-',    '-',    'S',    '-',    '-',    '-',  '-', '-', '-',    'S'  ));

CONSTANT udp_sedffsr : VitalStateTableType (1 TO 58, 1 TO 10) := ( 
--    NOTIFIER   D      CLK     RN       S      SI    SE   EN   Q(t)   Q(t+1)
     (  'X',    '-',    '-',    '-',    '-',    '-',  '-', '-', '-',    'X'  ),
     (  '-',    '-',    '-',    '0',    '1',    '-',  '-', '-', '-',    '0'  ), 
     (  '-',    '-',    '-',    '-',    '0',    '-',  '-', '-', '-',    '1'  ), 
     (  '-',    '-',    '/',    '-',    '1',    '0',  '1', '-', '-',    '0'  ),
     (  '-',    '-',    '/',    '1',    '-',    '1',  '1', '-', '-',    '1'  ), 
     (  '-',    '1',    '/',    '1',    '-',    '-',  '0', '1', '-',    '1'  ),
     (  '-',    '0',    '/',    '-',    '1',    '-',  '0', '1', '-',    '0'  ),
     (  '-',    '0',    '/',    '-',    '1',    '0',  '-', '1', '-',    '0'  ),
     (  '-',    '1',    '/',    '1',    '-',    '1',  '-', '1', '-',    '1'  ), 
     (  '-',    '-',    '-',    '1',    '-',    '-',  '0', '0', '1',    '1'  ), 
     (  '-',    '-',    '-',    '-',    '1',    '-',  '0', '0', '0',    '0'  ), 
     (  '-',    '-',    'X',    '1',    '-',    '1',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    'X',    '-',    '1',    '0',  '1', '-', '0',    '0'  ),
     (  '-',    '0',    'X',    '-',    '1',    '0',  '-', '-', '0',    '0'  ), 
     (  '-',    '1',    'X',    '1',    '-',    '1',  '-', '-', '1',    '1'  ), 
     (  '-',    '-',    'X',    '1',    '1',    '-',  '0', '0', '-',    'S'  ),
     (  '-',    '1',    'X',    '1',    '-',    '-',  '0', '-', '1',    '1'  ),-- no changes when in switches
     (  '-',    '1',    'X',    '-',    '1',    '-',  '0', '0', '0',    '0'  ),-- no changes when in switches
     (  '-',    '0',    'X',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),-- no changes when in switches
     (  '-',    '-',    '\',    '-',    '-',    '-',  '-', '-', '-',    'S'  ),-- no changes on falling clk edge
     (  '-',    '-',    '*',    '1',    '-',    '1',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '*',    '1',    '-',    '1',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '*',    '-',    '1',    '0',  '1', '-', '0',    '0'  ),
     (  '-',    '-',    '*',    '-',    '1',    '0',  '-', '0', '0',    '0'  ),
     (  '-',    '0',    '*',    '-',    '1',    '0',  '-', '-', '0',    '0'  ),
     (  '-',    '1',    '*',    '1',    '-',    '1',  '-', '-', '1',    '1'  ), 
     (  '-',    '-',    'S',    '1',    '-',    '-',  '*', '-', '1',    '1'  ),-- no changes when se switches
     (  '-',    '-',    'S',    '-',    '1',    '-',  '*', '-', '0',    '0'  ),-- no changes when se switches
     (  '-',    '-',    'S',    '-',    '1',    '*',  '-', '-', '0',    '0'  ),-- no changes when si switches
     (  '-',    '-',    'S',    '1',    '-',    '*',  '-', '-', '1',    '1'  ),-- no changes when si switches
     (  '-',    '*',    'S',    '1',    '-',    '-',  '-', '-', '1',    '1'  ),-- no changes when in switches
     (  '-',    '*',    'S',    '-',    '1',    '-',  '-', '-', '0',    '0'  ),-- no changes when in switches
     (  '-',    '*',    '-',    '1',    '-',    '1',  '-', '0', '1',    '1'  ),-- no changes when in switches
     (  '-',    '*',    '-',    '-',    '1',    '0',  '-', '0', '0',    '0'  ),-- no changes when in switches
     (  '-',    '-',    '-',    '1',    '-',    '1',  '*', '0', '1',    '1'  ),-- no changes when in switches
     (  '-',    '-',    '-',    '-',    '1',    '0',  '*', '0', '0',    '0'  ),-- no changes when in switches
     (  '-',    '-',    'S',    '1',    '-',    '-',  '-', '*', '1',    '1'  ),-- no changes when en switches
     (  '-',    '-',    'S',    '-',    '1',    '-',  '-', '*', '0',    '0'  ),-- no changes when en switches
     (  '-',    '-',    '*',    'B',    'B',    '-',  '0', '0', '-',    'S'  ), 
     (  '-',    '-',    '*',    'B',    'B',    '1',  '1', '-', '1',    '1'  ), 
     (  '-',    '-',    '*',    'B',    'B',    '0',  '1', '-', '0',    '0'  ), 
     (  '-',    '1',    '*',    'B',    'B',    '-',  '0', '1', '1',    '1'  ), 
     (  '-',    '0',    '*',    'B',    'B',    '-',  '0', '1', '0',    '0'  ), 
     (  '-',    '-',    '*',    '1',    '1',    '-',  '0', '0', '-',    'S'  ),
     (  '-',    '1',    '*',    '1',    '-',    '-',  '0', '-', '1',    '1'  ),-- reduce pessimism
     (  '-',    '0',    '*',    '-',    '1',    '-',  '0', '-', '0',    '0'  ),-- reduce pessimism
     (  '-',    '-',    '-',    '-',    '1',    '0',  '-', '0', '0',    '0'  ),-- reduce pessimism
     (  '-',    '-',    '-',    '1',    '-',    '1',  '-', '0', '1',    '1'  ),-- reduce pessimism
     (  '-',    '-',    '-',    '1',    '*',    '1',  '-', '0', '1',    '1'  ),
     (  '-',    '-',    '-',    '1',    '*',    '-',  '0', '0', '1',    '1'  ),
     (  '-',    '1',    '-',    '1',    '*',    '-',  '0', '1', '1',    '1'  ),
     (  '-',    '1',    '-',    '1',    '*',    '1',  '1', '-', '1',    '1'  ),
     (  '-',    '-',    '-',    '*',    '1',    '0',  '-', '0', '0',    '0'  ),
     (  '-',    '-',    '-',    '*',    '1',    '-',  '0', '0', '0',    '0'  ),
     (  '-',    '-',    '-',    '*',    '1',    '0',  '1', '-', '0',    '0'  ),
     (  '-',    '0',    '-',    '*',    '1',    '-',  '0', '1', '0',    '0'  ),
     (  '-',    '-',    'S',    '1',    '-',    '-',  '-', '-', '1',    '1'  ),
     (  '-',    '-',    'S',    '-',    '1',    '-',  '-', '-', '0',    '0'  ));

CONSTANT udp_pupd : VitalTruthTableType (1 TO 12, 1 TO 6) := (

    --  A       EN      PU      PD    data  control  
    
    (   '-',    '-',   '0',     '1',   'X',   'X' ),
    (   '-',    '-',   '0',     'X',   'X',   'X' ),
    (   '-',    '-',   'X',     '1',   'X',   'X' ),
    (   '-',    '-',   'X',     'X',   'X',   'X' ),

    (   '0',    '0',   '-',     '-',   '0',   '0' ),
    (   '0',    '1',   '-',     '-',   '0',   '1' ),
    (   '1',    '0',   '-',     '-',   '1',   '0' ),
    (   '1',    '1',   '-',     '-',   '1',   '1' ),
    (   '0',    'X',   '-',     '-',   '0',   'X' ),
    (   'X',    '0',   '-',     '-',   'X',   '0' ),
    (   '1',    'X',   '-',     '-',   '1',   'X' ),
    (   'X',    '1',   '-',     '-',   'X',   '1' ) );

CONSTANT udp_spupd : VitalTruthTableType (1 TO 16, 1 TO 7) := (
    --  S       A       EN      PU      PD    data  control  
    (   '-',   '-',    '-',   '0',     '1',   'X',   'X' ),
    (   '-',   '-',    '-',   '0',     'X',   'X',   'X' ),
    (   '-',   '-',    '-',   'X',     '1',   'X',   'X' ),
    (   '-',   '-',    '-',   'X',     'X',   'X',   'X' ),
    (   'X',   '0',    '0',   '-',     '-',   '0',   '0' ), -- added
    (   'X',   '1',    '0',   '-',     '-',   '1',   '0' ), -- added
    (   'X',   'X',    '0',   '-',     '-',   'X',   '0' ), -- added
    (   'X',   '-',    '-',   '-',     '-',   'X',   'X' ), -- added

    (   '-',   '0',    '0',   '-',     '-',   '0',   '0' ),
    (   '-',   '0',    '1',   '-',     '-',   '0',   '1' ),
    (   '-',   '1',    '0',   '-',     '-',   '1',   '0' ),
    (   '-',   '1',    '1',   '-',     '-',   '1',   '1' ),
    (   '-',   '0',    'X',   '-',     '-',   '0',   'X' ),
    (   '-',   'X',    '0',   '-',     '-',   'X',   '0' ),
    (   '-',   '1',    'X',   '-',     '-',   '1',   'X' ),
    (   '-',   'X',    '1',   '-',     '-',   'X',   '1' ) );

CONSTANT udp_sdpupd : VitalTruthTableType (1 TO 9, 1 TO 6) := (
    --  S      DLY     IN      PU      PD     out 
    (   'X',   '-',    '-',   '-',     '-',   'X' ),
    (   '-',   'X',    '-',   '-',     '-',   'X' ),
    (   '-',   '-',    '-',   '0',     '1',   'X' ),
    (   '-',   '-',    '-',   '0',     'X',   'X' ),
    (   '-',   '-',    '-',   'X',     '1',   'X' ),
    (   '-',   '-',    '-',   'X',     'X',   'X' ),
    (   '-',   '-',    '0',   '-',     '-',   '0' ),
    (   '-',   '-',    '1',   '-',     '-',   '1' ),
    (   '-',   '-',    'X',   '-',     '-',   'X' ));

CONSTANT udp_sdpupd_oe : VitalTruthTableType (1 TO 10, 1 TO 6) := (
    --  S      DLY     IN      PU      PD     out 
    (   '-',   '-',    '-',   '0',     '1',   'X' ),
    (   '-',   '-',    '-',   '0',     'X',   'X' ),
    (   '-',   '-',    '-',   'X',     '1',   'X' ),
    (   '-',   '-',    '-',   'X',     'X',   'X' ),
    (   'X',   '-',    '0',   '-',     '-',   '0' ),
    (   '-',   'X',    '-',   '-',     '-',   'X' ),
    (   'X',   '-',    '-',   '-',     '-',   'X' ),
    (   '-',   '-',    '0',   '-',     '-',   '0' ),
    (   '-',   '-',    '1',   '-',     '-',   '1' ),
    (   '-',   '-',    'X',   '-',     '-',   'X' ));

CONSTANT udp_dfflat : VitalStateTableType (1 TO 11, 1 TO 6) := (
--    NOTIFIER   D      CLK     CNTRL     Q(t)   Q(t+1)
    (   'X',    '-',    '-',    '-',      '-',    'X'  ),
    (   '-',    '0',    '-',    '1',      '-',    '0'  ),
    (   '-',    '1',    '-',    '1',      '-',    '1'  ),
    (   '-',    '1',    '/',    '0',      '-',    '1'  ),
    (   '-',    '0',    '/',    '0',      '-',    '0'  ),
    (   '-',    '1',    '*',    '0',      '1',    '1'  ),
    (   '-',    '0',    '*',    '0',      '0',    '0'  ),
    (   '-',    '-',    '\',    '0',      '-',    'S'  ),
    (   '-',    '-',    'B',    '0',      '-',    'S'  ),
    (   '-',    '*',    'B',    '0',      '-',    'S'  ),
    (   '-',    '-',    '-',    '/',      '-',    'S'  ));


end prim;

package body prim is

end prim;
--$Id: bmux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BENCX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_M2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_M2_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M2_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( 
            M2 : in std_ulogic := 'U';
            M1 : in std_ulogic := 'U';
            M0 : in std_ulogic := 'U';
            S : out std_ulogic;
            A : out std_ulogic;
            X2 : out std_ulogic);


     attribute VITAL_LEVEL0 of BENCX1 : entity is TRUE;
end BENCX1;

architecture behavioral of BENCX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL M2_ipd : std_ulogic := 'X';
     SIGNAL M1_ipd : std_ulogic := 'X';
     SIGNAL M0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( M2_ipd, M2, tipd_M2 );
          VitalWireDelay( M1_ipd, M1, tipd_M1 );
          VitalWireDelay( M0_ipd, M0, tipd_M0 );
END BLOCK;

VITALBehavior : PROCESS (M2_ipd, M1_ipd, M0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE S_zd : std_ulogic;
     VARIABLE A_zd : std_ulogic;
     VARIABLE X2_zd : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE A_GlitchData : VitalGlitchDataType;
     VARIABLE X2_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(M1_ipd);

          n1 := VitalINV(M0_ipd);

          n2 := VitalOR2(n0,n1);

          S_zd := VitalNAND2(M2_ipd,n2);
 
          n3 := VitalINV(M2_ipd);

          n4 := VitalOR2(M1_ipd, M0_ipd);

          A_zd := VitalNAND2(n3,n4);

          X2_zd := VitalXNOR2(M1_ipd, M0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_S,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_S,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_S,
                             TRUE)),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => A,
               OutSignalName => "A",
               OutTemp => A_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_A,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_A,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_A,
                             TRUE)),
               GlitchData => A_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => X2,
               OutSignalName => "X2",
               OutTemp => X2_zd,
               Paths => (
                      0 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_0,
                             (To_X01(M0_ipd) /= '1')),  
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_1,
                             (To_X01(M0_ipd) /= '0')),  
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_0,
                             (To_X01(M1_ipd) /= '1')),  
                      3 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_1,
                             (To_X01(M1_ipd) /= '0'))),  
               GlitchData => X2_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: bmux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BENCX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_M2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_M2_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M2_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( 
            M2 : in std_ulogic := 'U';
            M1 : in std_ulogic := 'U';
            M0 : in std_ulogic := 'U';
            S : out std_ulogic;
            A : out std_ulogic;
            X2 : out std_ulogic);


     attribute VITAL_LEVEL0 of BENCX2 : entity is TRUE;
end BENCX2;

architecture behavioral of BENCX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL M2_ipd : std_ulogic := 'X';
     SIGNAL M1_ipd : std_ulogic := 'X';
     SIGNAL M0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( M2_ipd, M2, tipd_M2 );
          VitalWireDelay( M1_ipd, M1, tipd_M1 );
          VitalWireDelay( M0_ipd, M0, tipd_M0 );
END BLOCK;

VITALBehavior : PROCESS (M2_ipd, M1_ipd, M0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE S_zd : std_ulogic;
     VARIABLE A_zd : std_ulogic;
     VARIABLE X2_zd : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE A_GlitchData : VitalGlitchDataType;
     VARIABLE X2_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(M1_ipd);

          n1 := VitalINV(M0_ipd);

          n2 := VitalOR2(n0,n1);

          S_zd := VitalNAND2(M2_ipd,n2);
 
          n3 := VitalINV(M2_ipd);

          n4 := VitalOR2(M1_ipd, M0_ipd);

          A_zd := VitalNAND2(n3,n4);

          X2_zd := VitalXNOR2(M1_ipd, M0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_S,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_S,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_S,
                             TRUE)),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => A,
               OutSignalName => "A",
               OutTemp => A_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_A,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_A,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_A,
                             TRUE)),
               GlitchData => A_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => X2,
               OutSignalName => "X2",
               OutTemp => X2_zd,
               Paths => (
                      0 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_0,
                             (To_X01(M0_ipd) /= '1')),  
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_1,
                             (To_X01(M0_ipd) /= '0')),  
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_0,
                             (To_X01(M1_ipd) /= '1')),  
                      3 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_1,
                             (To_X01(M1_ipd) /= '0'))),  
               GlitchData => X2_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: bmux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BENCX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_M2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_M2_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M2_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_A : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_X2_M1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_X2_M0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( 
            M2 : in std_ulogic := 'U';
            M1 : in std_ulogic := 'U';
            M0 : in std_ulogic := 'U';
            S : out std_ulogic;
            A : out std_ulogic;
            X2 : out std_ulogic);


     attribute VITAL_LEVEL0 of BENCX4 : entity is TRUE;
end BENCX4;

architecture behavioral of BENCX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL M2_ipd : std_ulogic := 'X';
     SIGNAL M1_ipd : std_ulogic := 'X';
     SIGNAL M0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( M2_ipd, M2, tipd_M2 );
          VitalWireDelay( M1_ipd, M1, tipd_M1 );
          VitalWireDelay( M0_ipd, M0, tipd_M0 );
END BLOCK;

VITALBehavior : PROCESS (M2_ipd, M1_ipd, M0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE S_zd : std_ulogic;
     VARIABLE A_zd : std_ulogic;
     VARIABLE X2_zd : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE A_GlitchData : VitalGlitchDataType;
     VARIABLE X2_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(M1_ipd);

          n1 := VitalINV(M0_ipd);

          n2 := VitalOR2(n0,n1);

          S_zd := VitalNAND2(M2_ipd,n2);
 
          n3 := VitalINV(M2_ipd);

          n4 := VitalOR2(M1_ipd, M0_ipd);

          A_zd := VitalNAND2(n3,n4);

          X2_zd := VitalXNOR2(M1_ipd, M0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_S,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_S,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_S,
                             TRUE)),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => A,
               OutSignalName => "A",
               OutTemp => A_zd,
               Paths => (
                      0 => ( M2_ipd'LAST_EVENT,
		             tpd_M2_A,
                             TRUE),
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_A,
                             TRUE),
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_A,
                             TRUE)),
               GlitchData => A_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => X2,
               OutSignalName => "X2",
               OutTemp => X2_zd,
               Paths => (
                      0 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_0,
                             (To_X01(M0_ipd) /= '1')),  
                      1 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_X2_M0_EQ_1,
                             (To_X01(M0_ipd) /= '0')),  
                      2 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_0,
                             (To_X01(M1_ipd) /= '1')),  
                      3 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_X2_M1_EQ_1,
                             (To_X01(M1_ipd) /= '0'))),  
               GlitchData => X2_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: bmux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BMXX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_M1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_M0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_X2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_A  : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_S  : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_PP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_PP_X2_EQ_1_AN_M0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_PP_X2_EQ_0_AN_M1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S_PP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S_PP_X2_EQ_1_AN_M0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S_PP_X2_EQ_0_AN_M1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_PP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_PP_X2_EQ_0_AN_A_EQ_1_AN_S_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M1_PP_X2_EQ_0_AN_A_EQ_0_AN_S_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_PP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_PP_X2_EQ_1_AN_A_EQ_1_AN_S_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_M0_PP_X2_EQ_1_AN_A_EQ_0_AN_S_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_X2_PP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_X2_PP_OP_M0_EQ_1_AN_A_EQ_1_AN_M1_EQ_0_AN_S_EQ_0_CP_OR_OP_M0_EQ_0_AN_S_EQ_1_AN_M1_EQ_1_AN_A_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_X2_PP_OP_M0_EQ_1_AN_A_EQ_0_AN_M1_EQ_0_AN_S_EQ_1_CP_OR_OP_M0_EQ_0_AN_S_EQ_0_AN_M1_EQ_1_AN_A_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( 
            X2 : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            S : in std_ulogic := 'U';
            M1 : in std_ulogic := 'U';
            M0 : in std_ulogic := 'U';
            PP : out std_ulogic);


     attribute VITAL_LEVEL0 of BMXX1 : entity is TRUE;
end BMXX1;

architecture behavioral of BMXX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL X2_ipd : std_ulogic := 'X';
     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL S_ipd : std_ulogic := 'X';
     SIGNAL M1_ipd : std_ulogic := 'X';
     SIGNAL M0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( X2_ipd, X2, tipd_X2 );
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( S_ipd, S, tipd_S );
          VitalWireDelay( M1_ipd, M1, tipd_M1 );
          VitalWireDelay( M0_ipd, M0, tipd_M0 );
END BLOCK;

VITALBehavior : PROCESS (X2_ipd, A_ipd, S_ipd, M1_ipd, M0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE PP_zd : std_ulogic;

     -- path delay section variables
     VARIABLE PP_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalTruthTable ( TruthTable => udp_bmx,
                                  DataIn => (X2_ipd, A_ipd, S_ipd, M1_ipd, M0_ipd));

          PP_zd := VitalBUF( n0 );

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => PP,
               OutSignalName => "PP",
               OutTemp => PP_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
		             tpd_A_PP_X2_EQ_1_AN_M0_EQ_1,
                             ((To_X01(X2_ipd) /= '0') and (To_X01(M0_ipd) /= '0'))),  
                      1 => ( A_ipd'LAST_EVENT,
		             tpd_A_PP_X2_EQ_0_AN_M1_EQ_1,
                             ((To_X01(X2_ipd) /= '1') and (To_X01(M1_ipd) /= '0'))),  
                      2 => ( S_ipd'LAST_EVENT,
		             tpd_S_PP_X2_EQ_1_AN_M0_EQ_0,
                             ((To_X01(X2_ipd) /= '0') and (To_X01(M0_ipd) /= '1'))),  
                      3 => ( S_ipd'LAST_EVENT,
		             tpd_S_PP_X2_EQ_0_AN_M1_EQ_0,
                             ((To_X01(X2_ipd) /= '1') and (To_X01(M1_ipd) /= '1'))),  
                      4 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_PP_X2_EQ_0_AN_A_EQ_1_AN_S_EQ_0,
                             ((To_X01(X2_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(S_ipd) /= '1'))),  
                      5 => ( M1_ipd'LAST_EVENT,
		             tpd_M1_PP_X2_EQ_0_AN_A_EQ_0_AN_S_EQ_1,
                             ((To_X01(X2_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(S_ipd) /= '0'))),  
                      6 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_PP_X2_EQ_1_AN_A_EQ_1_AN_S_EQ_0,
                             ((To_X01(X2_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(S_ipd) /= '1'))),  
                      7 => ( M0_ipd'LAST_EVENT,
		             tpd_M0_PP_X2_EQ_1_AN_A_EQ_0_AN_S_EQ_1,
                             ((To_X01(X2_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(S_ipd) /= '0'))),  
                      8 => ( X2_ipd'LAST_EVENT,
		             tpd_X2_PP_OP_M0_EQ_1_AN_A_EQ_1_AN_M1_EQ_0_AN_S_EQ_0_CP_OR_OP_M0_EQ_0_AN_S_EQ_1_AN_M1_EQ_1_AN_A_EQ_0_CP,
                             (((To_X01(M0_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(M1_ipd) /= '1') and (To_X01(S_ipd) /= '1')) or ((To_X01(M0_ipd) /= '1') and (To_X01(S_ipd) /= '0') and (To_X01(M1_ipd) /= '0') and (To_X01(A_ipd) /= '1')))),
                      9 => ( X2_ipd'LAST_EVENT,
		             tpd_X2_PP_OP_M0_EQ_1_AN_A_EQ_0_AN_M1_EQ_0_AN_S_EQ_1_CP_OR_OP_M0_EQ_0_AN_S_EQ_0_AN_M1_EQ_1_AN_A_EQ_1_CP,
                             (((To_X01(M0_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(M1_ipd) /= '1') and (To_X01(S_ipd) /= '0')) or ((To_X01(M0_ipd) /= '1') and (To_X01(S_ipd) /= '1') and (To_X01(M1_ipd) /= '0') and (To_X01(A_ipd) /= '0'))))),
               GlitchData => PP_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CMPR22X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of CMPR22X1 : entity is TRUE;
end CMPR22X1;

architecture behavioral of CMPR22X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,B_ipd);
 
          CO_zd := VitalAND2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: cmpr.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
use work.prim.all;

entity CMPR32X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( S : out std_ulogic;
            CO : out std_ulogic;
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of CMPR32X1 : entity is TRUE;
end CMPR32X1;

architecture behavioral of CMPR32X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,C_ipd);
 
          n0 := VitalAND2(A_ipd,B_ipd);

          n1 := VitalAND2(A_ipd,C_ipd);

          n2 := VitalAND2(B_ipd,C_ipd);

          CO_zd := VitalOR3(n0,n1,n2);



          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(C_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(C_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(C_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(C_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(C_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(C_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(C_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(C_ipd) /= '0'))),
                      8 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: cmpr.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
use work.prim.all;

entity CMPR42X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_ICI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_NT_OP_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_NT_OP_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_NT_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_NT_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( S : out std_ulogic;
            CO : out std_ulogic;
            ICO : out std_ulogic;
            ICI : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of CMPR42X1 : entity is TRUE;
end CMPR42X1;

architecture behavioral of CMPR42X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL ICI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( ICI_ipd, ICI, tipd_ICI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, ICI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE ICO_zd : std_ulogic;
     VARIABLE ISI : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;
     VARIABLE ICO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          ISI := VitalXOR3(A_ipd,B_ipd,C_ipd);

          n0 := VitalAND2(A_ipd,B_ipd);

          n1 := VitalAND2(A_ipd,C_ipd);

          n2 := VitalAND2(B_ipd,C_ipd);

          ICO_zd := VitalOR3(n0,n1,n2);

          S_zd := VitalXOR3(ISI,D_ipd,ICI_ipd);

          n3 := VitalAND2(ISI,D_ipd);

          n4 := VitalAND2(ISI,ICI_ipd);

          n5 := VitalAND2(D_ipd,ICI_ipd);

          CO_zd := VitalOR3(n3,n4,n5);
          


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1,
                             ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_NT_OP_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (NOT ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1,
                             ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_NT_OP_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))) or (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and (NOT ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))))),
                      5 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and (NOT((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))) or (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))))),

                      6 => ( D_ipd'LAST_EVENT,
                             tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and (To_X01(ICI_ipd) /= '0')) or ((NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0'))) and  (To_X01(ICI_ipd) /= '1')))),
                      7 => ( D_ipd'LAST_EVENT,
                             tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and (To_X01(ICI_ipd) /= '1')) or ((NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0'))) and  (To_X01(ICI_ipd) /= '0')))),
                      8 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_S_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1,
                             ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0'))),
                      9 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_CP,
                             (NOT(To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0')))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_NT_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_NT_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_CO_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      5 => ( C_ipd'LAST_EVENT,
                             tpd_C_CO_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      6 => ( D_ipd'LAST_EVENT,
                             tpd_D_CO,
                             TRUE ),
                      7 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => ICO,
               OutSignalName => "ICO",
               OutTemp => ICO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_ICO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_ICO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_ICO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_ICO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_ICO,
                             TRUE)),  
               GlitchData => ICO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: cmpr.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
use work.prim.all;

entity CMPR42X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_ICI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_NT_OP_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_NT_OP_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_ICO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_NT_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_NT_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_ICI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( S : out std_ulogic;
            CO : out std_ulogic;
            ICO : out std_ulogic;
            ICI : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of CMPR42X2 : entity is TRUE;
end CMPR42X2;

architecture behavioral of CMPR42X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL ICI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( ICI_ipd, ICI, tipd_ICI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, ICI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE ICO_zd : std_ulogic;
     VARIABLE ISI : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;
     VARIABLE ICO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          ISI := VitalXOR3(A_ipd,B_ipd,C_ipd);

          n0 := VitalAND2(A_ipd,B_ipd);

          n1 := VitalAND2(A_ipd,C_ipd);

          n2 := VitalAND2(B_ipd,C_ipd);

          ICO_zd := VitalOR3(n0,n1,n2);

          S_zd := VitalXOR3(ISI,D_ipd,ICI_ipd);

          n3 := VitalAND2(ISI,D_ipd);

          n4 := VitalAND2(ISI,ICI_ipd);

          n5 := VitalAND2(D_ipd,ICI_ipd);

          CO_zd := VitalOR3(n3,n4,n5);
          


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1,
                             ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_NT_OP_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (NOT ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1,
                             ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_NT_OP_A_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))) or (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and (NOT ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))))),
                      5 => ( C_ipd'LAST_EVENT,
                             tpd_C_S_OP_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_NT_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and (NOT((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))) or (NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0'))))),

                      6 => ( D_ipd'LAST_EVENT,
                             tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and (To_X01(ICI_ipd) /= '0')) or ((NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0'))) and  (To_X01(ICI_ipd) /= '1')))),
                      7 => ( D_ipd'LAST_EVENT,
                             tpd_D_S_OP_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_0_CP_OR_OP_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_CP_AN_ICI_EQ_1_CP,
                             ((((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and (To_X01(ICI_ipd) /= '1')) or ((NOT ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0'))) and  (To_X01(ICI_ipd) /= '0')))),
                      8 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_S_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1,
                             ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0'))),
                      9 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_C_EQ_1_XOB_D_EQ_1_CP,
                             (NOT(To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0') xor (To_X01(D_ipd) /= '0')))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_NT_OP_B_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(B_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_NT_OP_A_EQ_1_XOB_C_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(A_ipd) /= '0') xor (To_X01(C_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_CO_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      5 => ( C_ipd'LAST_EVENT,
                             tpd_C_CO_NT_OP_A_EQ_1_XOB_B_EQ_1_CP_AN_OP_D_EQ_1_XOB_ICI_EQ_1_CP,
                             (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')) and ((To_X01(D_ipd) /= '0') xor (To_X01(ICI_ipd) /= '0')))),
                      6 => ( D_ipd'LAST_EVENT,
                             tpd_D_CO,
                             TRUE ),
                      7 => ( ICI_ipd'LAST_EVENT,
                             tpd_ICI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => ICO,
               OutSignalName => "ICO",
               OutTemp => ICO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_ICO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_ICO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_ICO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_ICO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( C_ipd'LAST_EVENT,
                             tpd_C_ICO,
                             TRUE)),  
               GlitchData => ICO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFHCINX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CIN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_CIN_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CIN : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFHCINX2 : entity is TRUE;
end AFHCINX2;

architecture behavioral of AFHCINX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CIN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CIN_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CIN_ipd);

          n4 := VitalXOR2(A_ipd,B_ipd);
 
          S_zd := VitalXOR2(n4, n0);

          n1 := VitalAND2(A_ipd,B_ipd);

          n2 := VitalAND2(A_ipd,n0);

          n3 := VitalAND2(B_ipd,n0);
 
          CO_zd := VitalOR3(n3, n2, n1);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CIN_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CIN_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CIN_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CIN_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CIN_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CIN_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CIN_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CIN_ipd) /= '1'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CIN_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CIN_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CIN_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CIN_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CIN_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CIN_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CIN_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CIN_ipd) /= '1'))),
                      8 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFHCINX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CIN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_CIN_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CIN : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFHCINX4 : entity is TRUE;
end AFHCINX4;

architecture behavioral of AFHCINX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CIN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CIN_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CIN_ipd);

          n4 := VitalXOR2(A_ipd,B_ipd);
 
          S_zd := VitalXOR2(n4, n0);

          n1 := VitalAND2(A_ipd,B_ipd);

          n2 := VitalAND2(A_ipd,n0);

          n3 := VitalAND2(B_ipd,n0);
 
          CO_zd := VitalOR3(n3, n2, n1);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CIN_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CIN_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CIN_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CIN_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CIN_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CIN_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CIN_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CIN_ipd) /= '1'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CIN_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CIN_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CIN_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CIN_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CIN_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CIN_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CIN_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CIN_ipd) /= '1'))),
                      8 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFHCONX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CON : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFHCONX2 : entity is TRUE;
end AFHCONX2;

architecture behavioral of AFHCONX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CON_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CON_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n4 := VitalXOR2(A_ipd,B_ipd);
 
          S_zd := VitalXOR2(n4, CI_ipd);

          n1 := VitalAND2(A_ipd,B_ipd);

          n2 := VitalAND2(A_ipd,CI_ipd);

          n3 := VitalAND2(B_ipd,CI_ipd);
 
          CON_zd := VitalNOR3(n3, n2, n1);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CI_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CI_ipd) /= '1'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CI_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CI_ipd) /= '1'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CON,
               OutSignalName => "CON",
               OutTemp => CON_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CON_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CON_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CON,
                             TRUE )),
               GlitchData => CON_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFHCONX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CON_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CON : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFHCONX4 : entity is TRUE;
end AFHCONX4;

architecture behavioral of AFHCONX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CON_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CON_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n4 := VitalXOR2(A_ipd,B_ipd);
 
          S_zd := VitalXOR2(n4, CI_ipd);

          n1 := VitalAND2(A_ipd,B_ipd);

          n2 := VitalAND2(A_ipd,CI_ipd);

          n3 := VitalAND2(B_ipd,CI_ipd);
 
          CON_zd := VitalNOR3(n3, n2, n1);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CI_ipd) /= '0'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(CI_ipd) /= '1'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CI_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(CI_ipd) /= '1'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CON,
               OutSignalName => "CON",
               OutTemp => CON_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CON_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CON_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CON,
                             TRUE )),
               GlitchData => CON_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AHHCINX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CIN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            CIN : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AHHCINX2 : entity is TRUE;
end AHHCINX2;

architecture behavioral of AHHCINX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL CIN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, CIN_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CIN_ipd);

          S_zd := VitalXOR2(A_ipd,n0);

          CO_zd := VitalAND2(A_ipd,n0);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CIN_EQ_1,
                             (To_X01(CIN_ipd) /= '0')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CIN_EQ_0,
                             (To_X01(CIN_ipd) /= '1')),
                      2 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0')),
                      3 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AHHCINX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CIN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CIN_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CIN_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CIN_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            CIN : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AHHCINX4 : entity is TRUE;
end AHHCINX4;

architecture behavioral of AHHCINX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL CIN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( CIN_ipd, CIN, tipd_CIN );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, CIN_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CIN_ipd);

          S_zd := VitalXOR2(A_ipd,n0);

          CO_zd := VitalAND2(A_ipd,n0);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CIN_EQ_1,
                             (To_X01(CIN_ipd) /= '0')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CIN_EQ_0,
                             (To_X01(CIN_ipd) /= '1')),
                      2 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0')),
                      3 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( CIN_ipd'LAST_EVENT,
                             tpd_CIN_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AHHCONX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CON : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AHHCONX2 : entity is TRUE;
end AHHCONX2;

architecture behavioral of AHHCONX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CON_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CON_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,CI_ipd);

          CON_zd := VitalNAND2(A_ipd,CI_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CI_EQ_1,
                             (To_X01(CI_ipd) /= '0')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CI_EQ_0,
                             (To_X01(CI_ipd) /= '1')),
                      2 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0')),
                      3 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CON,
               OutSignalName => "CON",
               OutTemp => CON_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON,
                             TRUE ),
                      1 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CON,
                             TRUE )),
               GlitchData => CON_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AHHCONX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CON : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CON : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AHHCONX4 : entity is TRUE;
end AHHCONX4;

architecture behavioral of AHHCONX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CON_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CON_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,CI_ipd);

          CON_zd := VitalNAND2(A_ipd,CI_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CI_EQ_1,
                             (To_X01(CI_ipd) /= '0')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CI_EQ_0,
                             (To_X01(CI_ipd) /= '1')),
                      2 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0')),
                      3 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CON,
               OutSignalName => "CON",
               OutTemp => CON_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CON,
                             TRUE ),
                      1 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CON,
                             TRUE )),
               GlitchData => CON_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFCSHCINX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CS : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI0N : in std_ulogic := 'U';
            CI1N : in std_ulogic := 'U';
            CS : in std_ulogic := 'U';
            S : out std_ulogic;
            CO0 : out std_ulogic;
            CO1 : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFCSHCINX2 : entity is TRUE;
end AFCSHCINX2;

architecture behavioral of AFCSHCINX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI0N_ipd : std_ulogic := 'X';
     SIGNAL CI1N_ipd : std_ulogic := 'X';
     SIGNAL CS_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI0N_ipd, CI0N, tipd_CI0N );
          VitalWireDelay( CI1N_ipd, CI1N, tipd_CI1N );
          VitalWireDelay( CS_ipd, CS, tipd_CS );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI0N_ipd, CI1N_ipd, CS_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO0_zd : std_ulogic;
     VARIABLE CO1_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO0_GlitchData : VitalGlitchDataType;
     VARIABLE CO1_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CI0N_ipd);

          n1 := VitalINV(CI1N_ipd);

          n2 := VitalXOR3(A_ipd,B_ipd,n1);

          n3 := VitalAND2(CS_ipd,n2);

          n4 := VitalXOR3(A_ipd,B_ipd,n0);

          n5 := VitalINV(CS_ipd);

          n6 := VitalAND2(n5,n4);

          S_zd := VitalOR2(n6,n3);

          n7 := VitalAND2(A_ipd,B_ipd);

          n8 := VitalAND2(A_ipd,n0);

          n9 := VitalAND2(B_ipd,n0);
 
          CO0_zd := VitalOR3(n7, n8, n9);
          
          n10 := VitalAND2(A_ipd,B_ipd);

          n11 := VitalAND2(A_ipd,n1);

          n12 := VitalAND2(B_ipd,n1);
 
          CO1_zd := VitalOR3(n10, n11, n12);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1N_ipd) /= '0'))),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1N_ipd) /= '1'))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1N_ipd) /= '1'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1N_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0N_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0N_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0N_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0N_ipd) /= '0'))),
                      8 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1N_ipd) /= '0'))),
                      9 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1N_ipd) /= '1'))),
                      10 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1N_ipd) /= '1'))),
                      11 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1N_ipd) /= '0'))),
                      12 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0N_ipd) /= '0'))),
                      13 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0N_ipd) /= '1'))),
                      14 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0N_ipd) /= '1'))),
                      15 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0N_ipd) /= '0'))),
                      16 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      17 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      18 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      19 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      20 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1N_ipd) /= '1')) and (not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0N_ipd) /= '1'))))),
                      21 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP,
                             ((not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1N_ipd) /= '1'))) and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0N_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO0,
               OutSignalName => "CO0",
               OutTemp => CO0_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_CO0,
                             TRUE)),
               GlitchData => CO0_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO1,
               OutSignalName => "CO1",
               OutTemp => CO1_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_CO1,
                             TRUE)),
               GlitchData => CO1_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFCSHCINX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CS : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0N_CO0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1N_CO1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI0N : in std_ulogic := 'U';
            CI1N : in std_ulogic := 'U';
            CS : in std_ulogic := 'U';
            S : out std_ulogic;
            CO0 : out std_ulogic;
            CO1 : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFCSHCINX4 : entity is TRUE;
end AFCSHCINX4;

architecture behavioral of AFCSHCINX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI0N_ipd : std_ulogic := 'X';
     SIGNAL CI1N_ipd : std_ulogic := 'X';
     SIGNAL CS_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI0N_ipd, CI0N, tipd_CI0N );
          VitalWireDelay( CI1N_ipd, CI1N, tipd_CI1N );
          VitalWireDelay( CS_ipd, CS, tipd_CS );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI0N_ipd, CI1N_ipd, CS_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO0_zd : std_ulogic;
     VARIABLE CO1_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO0_GlitchData : VitalGlitchDataType;
     VARIABLE CO1_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalINV(CI0N_ipd);

          n1 := VitalINV(CI1N_ipd);

          n2 := VitalXOR3(A_ipd,B_ipd,n1);

          n3 := VitalAND2(CS_ipd,n2);

          n4 := VitalXOR3(A_ipd,B_ipd,n0);

          n5 := VitalINV(CS_ipd);

          n6 := VitalAND2(n5,n4);

          S_zd := VitalOR2(n6,n3);

          n7 := VitalAND2(A_ipd,B_ipd);

          n8 := VitalAND2(A_ipd,n0);

          n9 := VitalAND2(B_ipd,n0);
 
          CO0_zd := VitalOR3(n7, n8, n9);
          
          n10 := VitalAND2(A_ipd,B_ipd);

          n11 := VitalAND2(A_ipd,n1);

          n12 := VitalAND2(B_ipd,n1);
 
          CO1_zd := VitalOR3(n10, n11, n12);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1N_ipd) /= '0'))),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1N_ipd) /= '1'))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1N_ipd) /= '1'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1N_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0N_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0N_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0N_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0N_ipd) /= '0'))),
                      8 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1N_ipd) /= '0'))),
                      9 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1N_ipd) /= '1'))),
                      10 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1N_ipd) /= '1'))),
                      11 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1N_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1N_ipd) /= '0'))),
                      12 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0N_ipd) /= '0'))),
                      13 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0N_ipd) /= '1'))),
                      14 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0N_ipd) /= '1'))),
                      15 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0N_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0N_ipd) /= '0'))),
                      16 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      17 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      18 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      19 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      20 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1N_ipd) /= '1')) and (not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0N_ipd) /= '1'))))),
                      21 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1N_EQ_0_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0N_EQ_0_CP,
                             ((not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1N_ipd) /= '1'))) and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0N_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO0,
               OutSignalName => "CO0",
               OutTemp => CO0_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI0N_ipd'LAST_EVENT,
                             tpd_CI0N_CO0,
                             TRUE)),
               GlitchData => CO0_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO1,
               OutSignalName => "CO1",
               OutTemp => CO1_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI1N_ipd'LAST_EVENT,
                             tpd_CI1N_CO1,
                             TRUE)),
               GlitchData => CO1_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFCSHCONX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CS : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI0 : in std_ulogic := 'U';
            CI1 : in std_ulogic := 'U';
            CS : in std_ulogic := 'U';
            S : out std_ulogic;
            CO0N : out std_ulogic;
            CO1N : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFCSHCONX2 : entity is TRUE;
end AFCSHCONX2;

architecture behavioral of AFCSHCONX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI0_ipd : std_ulogic := 'X';
     SIGNAL CI1_ipd : std_ulogic := 'X';
     SIGNAL CS_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI0_ipd, CI0, tipd_CI0 );
          VitalWireDelay( CI1_ipd, CI1, tipd_CI1 );
          VitalWireDelay( CS_ipd, CS, tipd_CS );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI0_ipd, CI1_ipd, CS_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO0N_zd : std_ulogic;
     VARIABLE CO1N_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO0N_GlitchData : VitalGlitchDataType;
     VARIABLE CO1N_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n2 := VitalXOR3(A_ipd,B_ipd,CI1_ipd);

          n3 := VitalAND2(CS_ipd,n2);

          n4 := VitalXOR3(A_ipd,B_ipd,CI0_ipd);

          n5 := VitalINV(CS_ipd);

          n6 := VitalAND2(n5,n4);

          S_zd := VitalOR2(n6,n3);

          n7 := VitalAND2(A_ipd,B_ipd);

          n8 := VitalAND2(A_ipd,CI0_ipd);

          n9 := VitalAND2(B_ipd,CI0_ipd);
 
          CO0N_zd := VitalNOR3(n7, n8, n9);
          
          n10 := VitalAND2(A_ipd,B_ipd);

          n11 := VitalAND2(A_ipd,CI1_ipd);

          n12 := VitalAND2(B_ipd,CI1_ipd);
 
          CO1N_zd := VitalNOR3(n10, n11, n12);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1_ipd) /= '0'))),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1_ipd) /= '1'))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1_ipd) /= '1'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0_ipd) /= '0'))),
                      8 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1_ipd) /= '0'))),
                      9 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1_ipd) /= '1'))),
                      10 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1_ipd) /= '1'))),
                      11 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1_ipd) /= '0'))),
                      12 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0_ipd) /= '0'))),
                      13 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0_ipd) /= '1'))),
                      14 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0_ipd) /= '1'))),
                      15 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0_ipd) /= '0'))),
                      16 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      17 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      18 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      19 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      20 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1_ipd) /= '0')) and (not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0_ipd) /= '0'))))),
                      21 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP,
                             ((not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1_ipd) /= '0'))) and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0_ipd) /= '0'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO0N,
               OutSignalName => "CO0N",
               OutTemp => CO0N_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0N_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0N_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0N_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0N_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_CO0N,
                             TRUE)),
               GlitchData => CO0N_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO1N,
               OutSignalName => "CO1N",
               OutTemp => CO1N_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1N_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1N_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1N_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1N_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_CO1N,
                             TRUE)),
               GlitchData => CO1N_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AFCSHCONX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CS : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO0N_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO0N_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI0_CO0N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO1N_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO1N_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI1_CO1N : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI0 : in std_ulogic := 'U';
            CI1 : in std_ulogic := 'U';
            CS : in std_ulogic := 'U';
            S : out std_ulogic;
            CO0N : out std_ulogic;
            CO1N : out std_ulogic
            );

     attribute VITAL_LEVEL0 of AFCSHCONX4 : entity is TRUE;
end AFCSHCONX4;

architecture behavioral of AFCSHCONX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI0_ipd : std_ulogic := 'X';
     SIGNAL CI1_ipd : std_ulogic := 'X';
     SIGNAL CS_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI0_ipd, CI0, tipd_CI0 );
          VitalWireDelay( CI1_ipd, CI1, tipd_CI1 );
          VitalWireDelay( CS_ipd, CS, tipd_CS );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI0_ipd, CI1_ipd, CS_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO0N_zd : std_ulogic;
     VARIABLE CO1N_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO0N_GlitchData : VitalGlitchDataType;
     VARIABLE CO1N_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n2 := VitalXOR3(A_ipd,B_ipd,CI1_ipd);

          n3 := VitalAND2(CS_ipd,n2);

          n4 := VitalXOR3(A_ipd,B_ipd,CI0_ipd);

          n5 := VitalINV(CS_ipd);

          n6 := VitalAND2(n5,n4);

          S_zd := VitalOR2(n6,n3);

          n7 := VitalAND2(A_ipd,B_ipd);

          n8 := VitalAND2(A_ipd,CI0_ipd);

          n9 := VitalAND2(B_ipd,CI0_ipd);
 
          CO0N_zd := VitalNOR3(n7, n8, n9);
          
          n10 := VitalAND2(A_ipd,B_ipd);

          n11 := VitalAND2(A_ipd,CI1_ipd);

          n12 := VitalAND2(B_ipd,CI1_ipd);
 
          CO1N_zd := VitalNOR3(n10, n11, n12);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1_ipd) /= '0'))),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_0_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '1') and (To_X01(CI1_ipd) /= '1'))),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1_ipd) /= '1'))),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_1_AN_A_EQ_1_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(A_ipd) /= '0') and (To_X01(CI1_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0_ipd) /= '0'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_0_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '1') and (To_X01(CI0_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_CS_EQ_0_AN_A_EQ_1_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(A_ipd) /= '0') and (To_X01(CI0_ipd) /= '0'))),
                      8 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1_ipd) /= '0'))),
                      9 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_0_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '1') and (To_X01(CI1_ipd) /= '1'))),
                      10 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_0, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1_ipd) /= '1'))),
                      11 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_1_AN_B_EQ_1_AN_CI1_EQ_1, 
                             ((To_X01(CS_ipd) /= '0') and (To_X01(B_ipd) /= '0') and (To_X01(CI1_ipd) /= '0'))),
                      12 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0_ipd) /= '0'))),
                      13 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_0_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '1') and (To_X01(CI0_ipd) /= '1'))),
                      14 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_0, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0_ipd) /= '1'))),
                      15 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_CS_EQ_0_AN_B_EQ_1_AN_CI0_EQ_1, 
                             ((To_X01(CS_ipd) /= '1') and (To_X01(B_ipd) /= '0') and (To_X01(CI0_ipd) /= '0'))),
                      16 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_S_CS_EQ_0_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      17 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_S_CS_EQ_0_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '1') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      18 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_S_CS_EQ_1_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and (not ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0'))))),
                      19 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_S_CS_EQ_1_AN_OP_A_EQ_1_XOB_B_EQ_1_CP,
                             ((To_X01(CS_ipd) /= '0') and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0')))),
                      20 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP,
                             (((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1_ipd) /= '0')) and (not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0_ipd) /= '0'))))),
                      21 => ( CS_ipd'LAST_EVENT,
                             tpd_CS_S_NT_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI1_EQ_1_CP_AN_OP_A_EQ_1_XOB_B_EQ_1_XOB_CI0_EQ_1_CP,
                             ((not((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI1_ipd) /= '0'))) and ((To_X01(A_ipd) /= '0') xor (To_X01(B_ipd) /= '0') xor (To_X01(CI0_ipd) /= '0'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO0N,
               OutSignalName => "CO0N",
               OutTemp => CO0N_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0N_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO0N_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0N_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO0N_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI0_ipd'LAST_EVENT,
                             tpd_CI0_CO0N,
                             TRUE)),
               GlitchData => CO0N_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO1N,
               OutSignalName => "CO1N",
               OutTemp => CO1N_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1N_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO1N_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1N_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO1N_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI1_ipd'LAST_EVENT,
                             tpd_CI1_CO1N,
                             TRUE)),
               GlitchData => CO1N_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR3X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR3X2 : entity is TRUE;
end XNOR3X2;

architecture behavioral of XNOR3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd,C_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR3(A_ipd,B_ipd,C_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      8 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR3X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR3X4 : entity is TRUE;
end XNOR3X4;

architecture behavioral of XNOR3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd,C_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR3(A_ipd,B_ipd,C_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      8 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR3X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR3X2 : entity is TRUE;
end XOR3X2;

architecture behavioral of XOR3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd,C_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR3(A_ipd,B_ipd,C_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      8 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR3X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1_AN_C_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            C : in std_ulogic := 'U';
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR3X4 : entity is TRUE;
end XOR3X4;

architecture behavioral of XOR3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd,C_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR3(A_ipd,B_ipd,C_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_0,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1_AN_C_EQ_1,
                             ((To_X01(B_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '1'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(C_ipd) /= '0'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1_AN_C_EQ_1,
                             ((To_X01(A_ipd) /= '0') and (To_X01(C_ipd) /= '0'))),
                      8 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '1')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '0')))),
                      9 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0')) or ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1'))))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: rf.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
LIBRARY work;
USE work.prim.all;

entity RFRDX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_RB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RB_BRB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd)
              );

     port ( 
            RB : in std_ulogic := 'U';
            BRB : out std_ulogic
           );

     attribute VITAL_LEVEL0 of RFRDX1 : entity is TRUE;
end RFRDX1;

architecture behavioral of RFRDX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL io_wire : std_ulogic := 'X';
     CONSTANT ResultMapping : VitalResultMapType := ('W', 'W', 'L', 'H');
     SIGNAL RB_ipd : std_ulogic := 'X';


BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( RB_ipd, RB, tipd_RB );
END BLOCK;

VITALBehavior : PROCESS (RB_ipd)

     -- functionality section variables
     VARIABLE wwn : std_ulogic;
     VARIABLE BRB_zd : std_ulogic;

     -- path delay section variables
     VARIABLE BRB_GlitchData : VitalGlitchDataType;
     VARIABLE PrevData_udp_rfrd_n0 : std_logic_vector( 0 TO 1 );
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );

     VARIABLE n0 : std_ulogic := 'U';

     BEGIN
          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          VitalStateTable ( StateTable => udp_rfrd,
                           DataIn => ('1',RB_ipd),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_rfrd_n0 );

          n0 := n0_vec(1);
 
          BRB_zd := VitalBUF(n0);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => BRB,
               OutSignalName => "BRB",
               OutTemp => BRB_zd,
               Paths => (
                      0 => ( RB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_RB_BRB),
                             TRUE 
                            )),
               GlitchData => BRB_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: rf.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
LIBRARY work;
USE work.prim.all;

entity RFRDX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_RB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RB_BRB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd)
              );

     port ( 
            RB : in std_ulogic := 'U';
            BRB : out std_ulogic
           );

     attribute VITAL_LEVEL0 of RFRDX2 : entity is TRUE;
end RFRDX2;

architecture behavioral of RFRDX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL io_wire : std_ulogic := 'X';
     CONSTANT ResultMapping : VitalResultMapType := ('W', 'W', 'L', 'H');
     SIGNAL RB_ipd : std_ulogic := 'X';


BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( RB_ipd, RB, tipd_RB );
END BLOCK;

VITALBehavior : PROCESS (RB_ipd)

     -- functionality section variables
     VARIABLE wwn : std_ulogic;
     VARIABLE BRB_zd : std_ulogic;

     -- path delay section variables
     VARIABLE BRB_GlitchData : VitalGlitchDataType;
     VARIABLE PrevData_udp_rfrd_n0 : std_logic_vector( 0 TO 1 );
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );

     VARIABLE n0 : std_ulogic := 'U';

     BEGIN
          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          VitalStateTable ( StateTable => udp_rfrd,
                           DataIn => ('1',RB_ipd),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_rfrd_n0 );

          n0 := n0_vec(1);
 
          BRB_zd := VitalBUF(n0);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => BRB,
               OutSignalName => "BRB",
               OutTemp => BRB_zd,
               Paths => (
                      0 => ( RB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_RB_BRB),
                             TRUE 
                            )),
               GlitchData => BRB_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: rf.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
LIBRARY work;
USE work.prim.all;

entity RFRDX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_RB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RB_BRB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd)
              );

     port ( 
            RB : in std_ulogic := 'U';
            BRB : out std_ulogic
           );

     attribute VITAL_LEVEL0 of RFRDX4 : entity is TRUE;
end RFRDX4;

architecture behavioral of RFRDX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL io_wire : std_ulogic := 'X';
     CONSTANT ResultMapping : VitalResultMapType := ('W', 'W', 'L', 'H');
     SIGNAL RB_ipd : std_ulogic := 'X';


BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( RB_ipd, RB, tipd_RB );
END BLOCK;

VITALBehavior : PROCESS (RB_ipd)

     -- functionality section variables
     VARIABLE wwn : std_ulogic;
     VARIABLE BRB_zd : std_ulogic;

     -- path delay section variables
     VARIABLE BRB_GlitchData : VitalGlitchDataType;
     VARIABLE PrevData_udp_rfrd_n0 : std_logic_vector( 0 TO 1 );
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );

     VARIABLE n0 : std_ulogic := 'U';

     BEGIN
          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          VitalStateTable ( StateTable => udp_rfrd,
                           DataIn => ('1',RB_ipd),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_rfrd_n0 );

          n0 := n0_vec(1);
 
          BRB_zd := VitalBUF(n0);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => BRB,
               OutSignalName => "BRB",
               OutTemp => BRB_zd,
               Paths => (
                      0 => ( RB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_RB_BRB),
                             TRUE 
                            )),
               GlitchData => BRB_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: rf.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
LIBRARY work;
USE work.prim.all;

entity RF2R1WX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_WB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_WW : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_R1W : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_R2W : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tsetup_WB_WW_negedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_WB_WW_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_WB_WW_negedge_negedge : VitalDelayType := DefDummyHold;
               thold_WB_WW_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_WW_posedge : VitalDelayType := DefDummyWidth;
               tpd_WW_R1B : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_WW_R2B : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_WB_R1B : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_WB_R2B : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_R1W_R1B : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_R2W_R2B : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               TimingChecksOn : BOOLEAN := false
              );

     port ( 
            WB : in std_ulogic := 'U';
            WW : in std_ulogic := 'U';
            R1W : in std_ulogic := 'U';
            R2W : in std_ulogic := 'U';
            R1B : out std_ulogic;
            R2B : out std_ulogic
           );

     attribute VITAL_LEVEL0 of RF2R1WX2 : entity is TRUE;
end RF2R1WX2;

architecture behavioral of RF2R1WX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL WB_ipd : std_ulogic := 'X';
     SIGNAL WW_ipd : std_ulogic := 'X';
     SIGNAL R1W_ipd : std_ulogic := 'X';
     SIGNAL R2W_ipd : std_ulogic := 'X';


BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( WB_ipd, WB, tipd_WB );
          VitalWireDelay( WW_ipd, WW, tipd_WW );
          VitalWireDelay( R1W_ipd, R1W, tipd_R1W );
          VitalWireDelay( R2W_ipd, R2W, tipd_R2W );
END BLOCK;

VITALBehavior : PROCESS (WB_ipd, WW_ipd, R1W_ipd, R2W_ipd)

     -- timing checks section variables
     VARIABLE Tviol_WB_WW : std_ulogic := '0';
     VARIABLE TimeMarker_WB_WW : VitalTimingDataType;
     VARIABLE PWviol_WW_posedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_WW_posedge : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE wwn : std_ulogic;
     VARIABLE BRB_zd : std_ulogic;

     -- path delay section variables
     VARIABLE R1B_GlitchData : VitalGlitchDataType;
     VARIABLE R2B_GlitchData : VitalGlitchDataType;
     VARIABLE R1B_zd : std_ulogic;
     VARIABLE R2B_zd : std_ulogic;

     VARIABLE n0 : std_ulogic := 'U';
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE n1 : std_ulogic := 'U';
     VARIABLE n2 : std_ulogic := 'U';
     VARIABLE n3 : std_ulogic := 'U';
     VARIABLE n4 : std_ulogic := 'U';
     VARIABLE n5 : std_ulogic := 'U';
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlatrf_n0 : std_logic_vector( 0 TO 3 );
     VARIABLE PrevData_udp_tlatrf2_n0 : std_logic_vector( 0 TO 4 );

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => WB_ipd,
                   TestSignalName => "WB",
                   RefSignal      => WW_ipd,
                   RefSignalName  => "WW",
                   SetupHigh      => tsetup_WB_WW_posedge_negedge,
                   SetupLow       => tsetup_WB_WW_negedge_negedge,
                   HoldHigh       => thold_WB_WW_negedge_negedge,
                   HoldLow        => thold_WB_WW_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RF2R1WX2",
                   TimingData     => TimeMarker_WB_WW,
                   Violation      => Tviol_WB_WW,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => WW_ipd,
                   TestSignalName => "WW",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_WW_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_WW_posedge,
                   Violation      => PWviol_WW_posedge,
                   HeaderMsg      => InstancePath & "/RF2R1WX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_WB_WW OR 
                        PWviol_WW_posedge  
                       );
          n2 := VitalINV(WW_ipd); 

          n3 := VitalINV(R1W_ipd); 

          n4 := VitalINV(R2W_ipd); 

          VitalStateTable ( StateTable => udp_tlatrf,
                           DataIn => (NOTIFIER,WB_ipd,WW_ipd,n2),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlatrf_n0 );

          n0 := n0_vec(1);
          
          R1B_zd := VitalBUFIF1(n0, R1W_ipd);
 
          R2B_zd := VitalBUFIF1(n0, R2W_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => R1B,
               OutSignalName => "R1B",
               OutTemp => R1B_zd,
               Paths => (
                      0 => ( WW_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WW_R1B),
                             TRUE), 
                      1 => ( WB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WB_R1B),
                             TRUE), 
                      2 => ( R1W_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_R1W_R1B),
                             TRUE 
                            )),
               GlitchData => R1B_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01Z(
               OutSignal => R2B,
               OutSignalName => "R2B",
               OutTemp => R2B_zd,
               Paths => (
                      0 => ( WW_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WW_R2B),
                             TRUE), 
                      1 => ( WB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WB_R2B),
                             TRUE), 
                      2 => ( R2W_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_R2W_R2B),
                             TRUE 
                            )),
               GlitchData => R2B_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: rf.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
LIBRARY work;
USE work.prim.all;

entity RF1R1WX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_WB : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_WW : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_RW : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_RWN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tsetup_WB_WW_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_WB_WW_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_WB_WW_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_WB_WW_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_WW_posedge : VitalDelayType := DefDummyWidth;
               tpd_WW_RB : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_WB_RB : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_RW_RB : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_RWN_RB : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               TimingChecksOn : BOOLEAN := false
              );

     port ( 
            WB : in std_ulogic := 'U';
            WW : in std_ulogic := 'U';
            RW : in std_ulogic := 'U';
            RWN : in std_ulogic := 'U';
            RB : out std_ulogic
           );

     attribute VITAL_LEVEL0 of RF1R1WX2 : entity is TRUE;
end RF1R1WX2;

architecture behavioral of RF1R1WX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL WB_ipd : std_ulogic := 'X';
     SIGNAL WW_ipd : std_ulogic := 'X';
     SIGNAL RW_ipd : std_ulogic := 'X';
     SIGNAL RWN_ipd : std_ulogic := 'X';


BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( WB_ipd, WB, tipd_WB );
          VitalWireDelay( WW_ipd, WW, tipd_WW );
          VitalWireDelay( RW_ipd, RW, tipd_RW );
          VitalWireDelay( RWN_ipd, RWN, tipd_RWN );
END BLOCK;

VITALBehavior : PROCESS (WB_ipd, WW_ipd, RW_ipd, RWN_ipd)

     -- timing checks section variables
     VARIABLE Tviol_WB_WW : std_ulogic := '0';
     VARIABLE TimeMarker_WB_WW : VitalTimingDataType;
     VARIABLE PWviol_WW_posedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_WW_posedge : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE wwn : std_ulogic;
     VARIABLE BRB_zd : std_ulogic;

     -- path delay section variables
     VARIABLE RB_GlitchData : VitalGlitchDataType;
     VARIABLE RB_zd : std_ulogic;

     VARIABLE n0 : std_ulogic := 'U';
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE n1 : std_ulogic := 'U';
     VARIABLE n2 : std_ulogic := 'U';
     VARIABLE n3 : std_ulogic := 'U';
     VARIABLE n4 : std_ulogic := 'U';
     VARIABLE n5 : std_ulogic := 'U';
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlatrf_n0 : std_logic_vector( 0 TO 3 );
     VARIABLE PrevData_udp_tlatrf2_n0 : std_logic_vector( 0 TO 4 );

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => WB_ipd,
                   TestSignalName => "WB",
                   RefSignal      => WW_ipd,
                   RefSignalName  => "WW",
                   SetupHigh      => tsetup_WB_WW_posedge_negedge,
                   SetupLow       => tsetup_WB_WW_negedge_negedge,
                   HoldHigh       => thold_WB_WW_negedge_negedge,
                   HoldLow        => thold_WB_WW_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RF1R1WX2",
                   TimingData     => TimeMarker_WB_WW,
                   Violation      => Tviol_WB_WW,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => WW_ipd,
                   TestSignalName => "WW",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_WW_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_WW_posedge,
                   Violation      => PWviol_WW_posedge,
                   HeaderMsg      => InstancePath & "/RF1R1WX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_WB_WW OR 
                        PWviol_WW_posedge 
                       );

          wwn := VitalINV(WW_ipd);

          VitalStateTable ( StateTable => udp_tlatrf,
                           DataIn => (NOTIFIER,WB_ipd,WW_ipd,wwn),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlatrf_n0 );

          n0 := n0_vec(1);
          
          n1 := VitalTruthTable ( TruthTable => udp_outrf,
                                  DataIn => (n0,RW_ipd,RWN_ipd));

          RB_zd := VitalBUFIF1(n0, n1);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => RB,
               OutSignalName => "RB",
               OutTemp => RB_zd,
               Paths => (
                      0 => ( WW_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WW_RB),
                             TRUE), 
                      1 => ( WB_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_WB_RB),
                             TRUE), 
                      2 => ( RW_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_RW_RB),
                             TRUE), 
                      3 => ( RWN_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_RWN_RB),
                             TRUE 
                            )),
               GlitchData => RB_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;
--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFHX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFHX1 : entity is TRUE;
end ADDFHX1;

architecture behavioral of ADDFHX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFHX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFHX2 : entity is TRUE;
end ADDFHX2;

architecture behavioral of ADDFHX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFHX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFHX4 : entity is TRUE;
end ADDFHX4;

architecture behavioral of ADDFHX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFHXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFHXL : entity is TRUE;
end ADDFHXL;

architecture behavioral of ADDFHXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFX1 : entity is TRUE;
end ADDFX1;

architecture behavioral of ADDFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFX2 : entity is TRUE;
end ADDFX2;

architecture behavioral of ADDFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFX4 : entity is TRUE;
end ADDFX4;

architecture behavioral of ADDFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDFXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_CO_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1_AN_CI_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CI_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            CI : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDFXL : entity is TRUE;
end ADDFXL;

architecture behavioral of ADDFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL CI_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( CI_ipd, CI, tipd_CI );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, CI_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE a_and_b : std_ulogic;
     VARIABLE a_and_ci : std_ulogic;
     VARIABLE b_and_ci : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR3(A_ipd,B_ipd,CI_ipd);

          a_and_b := VitalAND2(A_ipd,B_ipd);

          a_and_ci := VitalAND2(A_ipd,CI_ipd);

          b_and_ci := VitalAND2(B_ipd,CI_ipd);

          CO_zd := VitalOR3(a_and_b,a_and_ci,b_and_ci);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      2 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_0,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      3 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1_AN_CI_EQ_1,
                             ((To_X01(B_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      4 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '1'))),
                      5 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '1') AND (To_X01(CI_ipd) /= '0'))),
                      6 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_0,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '1'))),
                      7 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1_AN_CI_EQ_1,
                             ((To_X01(A_ipd) /= '0') AND (To_X01(CI_ipd) /= '0'))),
                      8 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_1_CP_OR_OP_A_EQ_1_AN_B_EQ_0_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '1')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '0')))),
                      9 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_S_OP_A_EQ_0_AN_B_EQ_0_CP_OR_OP_A_EQ_1_AN_B_EQ_1_CP,
                             (((To_X01(B_ipd) /= '0') AND (To_X01(A_ipd) /= '0')) OR ((To_X01(B_ipd) /= '1') AND (To_X01(A_ipd) /= '1'))))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_0,
                             (To_X01(B_ipd) /= '1') ),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO_B_EQ_1,
                             (To_X01(B_ipd) /= '0') ),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_0,
                             (To_X01(A_ipd) /= '1') ),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO_A_EQ_1,
                             (To_X01(A_ipd) /= '0') ),
                      4 => ( CI_ipd'LAST_EVENT,
                             tpd_CI_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDHX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDHX1 : entity is TRUE;
end ADDHX1;

architecture behavioral of ADDHX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,B_ipd);
 
          CO_zd := VitalAND2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDHX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDHX2 : entity is TRUE;
end ADDHX2;

architecture behavioral of ADDHX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,B_ipd);
 
          CO_zd := VitalAND2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDHX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDHX4 : entity is TRUE;
end ADDHX4;

architecture behavioral of ADDHX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,B_ipd);
 
          CO_zd := VitalAND2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: add.genpp,v 1.3 2001/08/23 18:37:12 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity ADDHXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_S_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_S_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_CO : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S : out std_ulogic;
            CO : out std_ulogic
            );

     attribute VITAL_LEVEL0 of ADDHXL : entity is TRUE;
end ADDHXL;

architecture behavioral of ADDHXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE S_zd : std_ulogic;
     VARIABLE CO_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE n2 : std_ulogic;
     VARIABLE n3 : std_ulogic;
     VARIABLE n4 : std_ulogic;
     VARIABLE n5 : std_ulogic;
     VARIABLE n6 : std_ulogic;
     VARIABLE n7 : std_ulogic;
     VARIABLE n8 : std_ulogic;
     VARIABLE n9 : std_ulogic;
     VARIABLE n10 : std_ulogic;
     VARIABLE n11 : std_ulogic;
     VARIABLE n12 : std_ulogic;
     VARIABLE n13 : std_ulogic;
     VARIABLE n14 : std_ulogic;

     -- path delay section variables
     VARIABLE S_GlitchData : VitalGlitchDataType;
     VARIABLE CO_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          S_zd := VitalXOR2(A_ipd,B_ipd);
 
          CO_zd := VitalAND2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => S,
               OutSignalName => "S",
               OutTemp => S_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_S_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_S_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => S_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => CO,
               OutSignalName => "CO",
               OutTemp => CO_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_CO,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_CO,
                             TRUE )),
               GlitchData => CO_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


END PROCESS;
end behavioral;

--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND2X1 : entity is TRUE;
end AND2X1;

architecture behavioral of AND2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND2X2 : entity is TRUE;
end AND2X2;

architecture behavioral of AND2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND2X4 : entity is TRUE;
end AND2X4;

architecture behavioral of AND2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND2XL : entity is TRUE;
end AND2XL;

architecture behavioral of AND2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND3X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND3X1 : entity is TRUE;
end AND3X1;

architecture behavioral of AND3X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND3X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND3X2 : entity is TRUE;
end AND3X2;

architecture behavioral of AND3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND3X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND3X4 : entity is TRUE;
end AND3X4;

architecture behavioral of AND3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND3XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND3XL : entity is TRUE;
end AND3XL;

architecture behavioral of AND3XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND4X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND4X1 : entity is TRUE;
end AND4X1;

architecture behavioral of AND4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND4X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND4X2 : entity is TRUE;
end AND4X2;

architecture behavioral of AND4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND4X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND4X4 : entity is TRUE;
end AND4X4;

architecture behavioral of AND4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AND4XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AND4XL : entity is TRUE;
end AND4XL;

architecture behavioral of AND4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI211X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI211X1 : entity is TRUE;
end AOI211X1;

architecture behavioral of AOI211X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI211X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI211X2 : entity is TRUE;
end AOI211X2;

architecture behavioral of AOI211X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI211X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI211X4 : entity is TRUE;
end AOI211X4;

architecture behavioral of AOI211X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI211XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI211XL : entity is TRUE;
end AOI211XL;

architecture behavioral of AOI211XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI21X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI21X1 : entity is TRUE;
end AOI21X1;

architecture behavioral of AOI21X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI21X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI21X2 : entity is TRUE;
end AOI21X2;

architecture behavioral of AOI21X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI21X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI21X4 : entity is TRUE;
end AOI21X4;

architecture behavioral of AOI21X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI21XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI21XL : entity is TRUE;
end AOI21XL;

architecture behavioral of AOI21XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI221X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI221X1 : entity is TRUE;
end AOI221X1;

architecture behavioral of AOI221X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI221X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI221X2 : entity is TRUE;
end AOI221X2;

architecture behavioral of AOI221X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI221X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI221X4 : entity is TRUE;
end AOI221X4;

architecture behavioral of AOI221X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI221XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI221XL : entity is TRUE;
end AOI221XL;

architecture behavioral of AOI221XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI222X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI222X1 : entity is TRUE;
end AOI222X1;

architecture behavioral of AOI222X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          outC := VitalAND2(C0_ipd, C1_ipd);

          Y_zd := VitalNOR3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI222X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI222X2 : entity is TRUE;
end AOI222X2;

architecture behavioral of AOI222X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          outC := VitalAND2(C0_ipd, C1_ipd);

          Y_zd := VitalNOR3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI222X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI222X4 : entity is TRUE;
end AOI222X4;

architecture behavioral of AOI222X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          outC := VitalAND2(C0_ipd, C1_ipd);

          Y_zd := VitalNOR3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI222XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI222XL : entity is TRUE;
end AOI222XL;

architecture behavioral of AOI222XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          outC := VitalAND2(C0_ipd, C1_ipd);

          Y_zd := VitalNOR3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI22X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI22X1 : entity is TRUE;
end AOI22X1;

architecture behavioral of AOI22X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI22X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI22X2 : entity is TRUE;
end AOI22X2;

architecture behavioral of AOI22X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI22X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI22X4 : entity is TRUE;
end AOI22X4;

architecture behavioral of AOI22X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI22XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI22XL : entity is TRUE;
end AOI22XL;

architecture behavioral of AOI22XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND2(A0_ipd, A1_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB1X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB1X1 : entity is TRUE;
end AOI2BB1X1;

architecture behavioral of AOI2BB1X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB1X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB1X2 : entity is TRUE;
end AOI2BB1X2;

architecture behavioral of AOI2BB1X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB1X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB1X4 : entity is TRUE;
end AOI2BB1X4;

architecture behavioral of AOI2BB1X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB1XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB1XL : entity is TRUE;
end AOI2BB1XL;

architecture behavioral of AOI2BB1XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB2X1 : entity is TRUE;
end AOI2BB2X1;

architecture behavioral of AOI2BB2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB2X2 : entity is TRUE;
end AOI2BB2X2;

architecture behavioral of AOI2BB2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB2X4 : entity is TRUE;
end AOI2BB2X4;

architecture behavioral of AOI2BB2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI2BB2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI2BB2XL : entity is TRUE;
end AOI2BB2XL;

architecture behavioral of AOI2BB2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalAND2(A0X_ipd, A1X_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI31X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI31X1 : entity is TRUE;
end AOI31X1;

architecture behavioral of AOI31X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI31X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI31X2 : entity is TRUE;
end AOI31X2;

architecture behavioral of AOI31X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI31X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI31X4 : entity is TRUE;
end AOI31X4;

architecture behavioral of AOI31X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI31XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI31XL : entity is TRUE;
end AOI31XL;

architecture behavioral of AOI31XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNOR2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI32X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI32X1 : entity is TRUE;
end AOI32X1;

architecture behavioral of AOI32X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI32X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI32X2 : entity is TRUE;
end AOI32X2;

architecture behavioral of AOI32X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI32X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI32X4 : entity is TRUE;
end AOI32X4;

architecture behavioral of AOI32X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI32XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI32XL : entity is TRUE;
end AOI32XL;

architecture behavioral of AOI32XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND2(B0_ipd, B1_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI33X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI33X1 : entity is TRUE;
end AOI33X1;

architecture behavioral of AOI33X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI33X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI33X2 : entity is TRUE;
end AOI33X2;

architecture behavioral of AOI33X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI33X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI33X4 : entity is TRUE;
end AOI33X4;

architecture behavioral of AOI33X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity AOI33XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of AOI33XL : entity is TRUE;
end AOI33XL;

architecture behavioral of AOI33XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalAND3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalAND3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNOR2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX12 : entity is TRUE;
end BUFX12;

architecture behavioral of BUFX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX16 : entity is TRUE;
end BUFX16;

architecture behavioral of BUFX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX1 : entity is TRUE;
end BUFX1;

architecture behavioral of BUFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX20 : entity is TRUE;
end BUFX20;

architecture behavioral of BUFX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX2 : entity is TRUE;
end BUFX2;

architecture behavioral of BUFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX3 : entity is TRUE;
end BUFX3;

architecture behavioral of BUFX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX4 : entity is TRUE;
end BUFX4;

architecture behavioral of BUFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFX8 : entity is TRUE;
end BUFX8;

architecture behavioral of BUFX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity BUFXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of BUFXL : entity is TRUE;
end BUFXL;

architecture behavioral of BUFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX12 : entity is TRUE;
end CLKBUFX12;

architecture behavioral of CLKBUFX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX16 : entity is TRUE;
end CLKBUFX16;

architecture behavioral of CLKBUFX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX1 : entity is TRUE;
end CLKBUFX1;

architecture behavioral of CLKBUFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX20 : entity is TRUE;
end CLKBUFX20;

architecture behavioral of CLKBUFX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX2 : entity is TRUE;
end CLKBUFX2;

architecture behavioral of CLKBUFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX3 : entity is TRUE;
end CLKBUFX3;

architecture behavioral of CLKBUFX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX4 : entity is TRUE;
end CLKBUFX4;

architecture behavioral of CLKBUFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFX8 : entity is TRUE;
end CLKBUFX8;

architecture behavioral of CLKBUFX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKBUFXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKBUFXL : entity is TRUE;
end CLKBUFXL;

architecture behavioral of CLKBUFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX12 : entity is TRUE;
end CLKINVX12;

architecture behavioral of CLKINVX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX16 : entity is TRUE;
end CLKINVX16;

architecture behavioral of CLKINVX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX1 : entity is TRUE;
end CLKINVX1;

architecture behavioral of CLKINVX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX20 : entity is TRUE;
end CLKINVX20;

architecture behavioral of CLKINVX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX2 : entity is TRUE;
end CLKINVX2;

architecture behavioral of CLKINVX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX3 : entity is TRUE;
end CLKINVX3;

architecture behavioral of CLKINVX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX4 : entity is TRUE;
end CLKINVX4;

architecture behavioral of CLKINVX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVX8 : entity is TRUE;
end CLKINVX8;

architecture behavioral of CLKINVX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity CLKINVXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of CLKINVXL : entity is TRUE;
end CLKINVXL;

architecture behavioral of CLKINVXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFX1 : entity is TRUE;
end DFFX1;

architecture behavioral of DFFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFX2 : entity is TRUE;
end DFFX2;

architecture behavioral of DFFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFX4 : entity is TRUE;
end DFFX4;

architecture behavioral of DFFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFXL : entity is TRUE;
end DFFXL;

architecture behavioral of DFFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFHQX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFHQX1 : entity is TRUE;
end DFFHQX1;

architecture behavioral of DFFHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFHQX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFHQX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFHQX2 : entity is TRUE;
end DFFHQX2;

architecture behavioral of DFFHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFHQX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFHQX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFHQX4 : entity is TRUE;
end DFFHQX4;

architecture behavioral of DFFHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFHQX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFHQXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFHQXL : entity is TRUE;
end DFFHQXL;

architecture behavioral of DFFHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFHQXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNX1 : entity is TRUE;
end DFFNX1;

architecture behavioral of DFFNX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNX2 : entity is TRUE;
end DFFNX2;

architecture behavioral of DFFNX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNX4 : entity is TRUE;
end DFFNX4;

architecture behavioral of DFFNX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNXL : entity is TRUE;
end DFFNXL;

architecture behavioral of DFFNXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNRX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNRX1 : entity is TRUE;
end DFFNRX1;

architecture behavioral of DFFNRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX1",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNRX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNRX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNRX2 : entity is TRUE;
end DFFNRX2;

architecture behavioral of DFFNRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX2",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNRX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNRX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNRX4 : entity is TRUE;
end DFFNRX4;

architecture behavioral of DFFNRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX4",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNRX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNRXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNRXL : entity is TRUE;
end DFFNRXL;

architecture behavioral of DFFNRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRXL",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNRXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNRXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSX1 : entity is TRUE;
end DFFNSX1;

architecture behavioral of DFFNSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX1",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSX2 : entity is TRUE;
end DFFNSX2;

architecture behavioral of DFFNSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX2",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSX4 : entity is TRUE;
end DFFNSX4;

architecture behavioral of DFFNSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX4",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSXL : entity is TRUE;
end DFFNSXL;

architecture behavioral of DFFNSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSXL",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSRX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSRX1 : entity is TRUE;
end DFFNSRX1;

architecture behavioral of DFFNSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSRX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSRX2 : entity is TRUE;
end DFFNSRX2;

architecture behavioral of DFFNSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSRX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSRX4 : entity is TRUE;
end DFFNSRX4;

architecture behavioral of DFFNSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFNSRXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFNSRXL : entity is TRUE;
end DFFNSRXL;

architecture behavioral of DFFNSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   TimingData     => TimeMarker_RN_CKN,
                   Violation      => Tviol_RN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CKN_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   TimingData     => TimeMarker_SN_CKN,
                   Violation      => Tviol_SN_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRX1 : entity is TRUE;
end DFFRX1;

architecture behavioral of DFFRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRX2 : entity is TRUE;
end DFFRX2;

architecture behavioral of DFFRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRX4 : entity is TRUE;
end DFFRX4;

architecture behavioral of DFFRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRXL : entity is TRUE;
end DFFRXL;

architecture behavioral of DFFRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRHQX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRHQX1 : entity is TRUE;
end DFFRHQX1;

architecture behavioral of DFFRHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRHQX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRHQX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRHQX2 : entity is TRUE;
end DFFRHQX2;

architecture behavioral of DFFRHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRHQX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRHQX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRHQX4 : entity is TRUE;
end DFFRHQX4;

architecture behavioral of DFFRHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRHQX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFRHQXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFRHQXL : entity is TRUE;
end DFFRHQXL;

architecture behavioral of DFFRHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFRHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFRHQXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSX1 : entity is TRUE;
end DFFSX1;

architecture behavioral of DFFSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSX2 : entity is TRUE;
end DFFSX2;

architecture behavioral of DFFSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSX4 : entity is TRUE;
end DFFSX4;

architecture behavioral of DFFSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSXL : entity is TRUE;
end DFFSXL;

architecture behavioral of DFFSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSHQX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSHQX1 : entity is TRUE;
end DFFSHQX1;

architecture behavioral of DFFSHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSHQX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSHQX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSHQX2 : entity is TRUE;
end DFFSHQX2;

architecture behavioral of DFFSHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSHQX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSHQX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSHQX4 : entity is TRUE;
end DFFSHQX4;

architecture behavioral of DFFSHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSHQX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSHQXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSHQXL : entity is TRUE;
end DFFSHQXL;

architecture behavioral of DFFSHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSHQXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRX1 : entity is TRUE;
end DFFSRX1;

architecture behavioral of DFFSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRX2 : entity is TRUE;
end DFFSRX2;

architecture behavioral of DFFSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRX4 : entity is TRUE;
end DFFSRX4;

architecture behavioral of DFFSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRXL : entity is TRUE;
end DFFSRXL;

architecture behavioral of DFFSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRHQX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRHQX1 : entity is TRUE;
end DFFSRHQX1;

architecture behavioral of DFFSRHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRHQX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRHQX2 : entity is TRUE;
end DFFSRHQX2;

architecture behavioral of DFFSRHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRHQX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRHQX4 : entity is TRUE;
end DFFSRHQX4;

architecture behavioral of DFFSRHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFSRHQXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFSRHQXL : entity is TRUE;
end DFFSRHQXL;

architecture behavioral of DFFSRHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/DFFSRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_RN OR 
                        Tviol_RN_SN OR 
                        Tviol_D_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,D_dly,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(flag) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFTRX1 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFTRX1 : entity is TRUE;
end DFFTRX1;

architecture behavioral of DFFTRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE E : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => To_X01(D_dly) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFTRX1",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          E := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFTRX2 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFTRX2 : entity is TRUE;
end DFFTRX2;

architecture behavioral of DFFTRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE E : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => To_X01(D_dly) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFTRX2",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          E := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFTRX4 is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFTRX4 : entity is TRUE;
end DFFTRX4;

architecture behavioral of DFFTRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE E : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => To_X01(D_dly) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFTRX4",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          E := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: dff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DFFTRXL is

     generic ( 
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               ticd_CK : VitalDelayType := DefDummyIcd;
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of DFFTRXL : entity is TRUE;
end DFFTRXL;

architecture behavioral of DFFTRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;

     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE intclk : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE E : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE QN_GlitchData : VitalGlitchDataType;
     VARIABLE QN_zd : std_ulogic;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => To_X01(D_dly) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/DFFTRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/DFFTRXL",
                   CheckEnabled   => ( To_X01(flag) ) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          E := '1';

          intclk := VitalBUF(CK_dly);

 
          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );

          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );
 
          flag := VitalAND2(SNx_dly,RNx_dly);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DLY1X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of DLY1X1 : entity is TRUE;
end DLY1X1;

architecture behavioral of DLY1X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DLY2X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of DLY2X1 : entity is TRUE;
end DLY2X1;

architecture behavioral of DLY2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DLY3X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of DLY3X1 : entity is TRUE;
end DLY3X1;

architecture behavioral of DLY3X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity DLY4X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of DLY4X1 : entity is TRUE;
end DLY4X1;

architecture behavioral of DLY4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUF(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFX1 : entity is TRUE;
end EDFFX1;

architecture behavioral of EDFFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX1",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFX2 : entity is TRUE;
end EDFFX2;

architecture behavioral of EDFFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX2",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFX4 : entity is TRUE;
end EDFFX4;

architecture behavioral of EDFFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFX4",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFXL : entity is TRUE;
end EDFFXL;

architecture behavioral of EDFFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFXL",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFTRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFTRX1 : entity is TRUE;
end EDFFTRX1;

architecture behavioral of EDFFTRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX1",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFTRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFTRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFTRX2 : entity is TRUE;
end EDFFTRX2;

architecture behavioral of EDFFTRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX2",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFTRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFTRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFTRX4 : entity is TRUE;
end EDFFTRX4;

architecture behavioral of EDFFTRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX4",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFTRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity EDFFTRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of EDFFTRXL : entity is TRUE;
end EDFFTRXL;

architecture behavioral of EDFFTRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE SIx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_edfft_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRXL",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/EDFFTRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/EDFFTRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_edfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_edfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := '1';

          SIx_dly := VitalBUF( D_dly);

          DxorSI := VitalXOR2(D_dly, SIx_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

--LIBRARY IEEE;
--USE IEEE.Std_logic_1164.all;
--USE IEEE.VITAL_Timing.all;
--USE IEEE.VITAL_Primitives.all;
--USE work.prim.all;
--
--entity HOLDX1 is
--
--     generic ( 
--               XOn    : BOOLEAN := DefCombSpikeXOn;
--               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
--               InstancePath : STRING := "*";
--               tipd_Y : VitalDelayType01 := (DefDummyIpd, DefDummyIpd)
--              );
--
--     port ( 
--            Y : inout std_ulogic
--           );
--
--     attribute VITAL_LEVEL0 of HOLDX1 : entity is TRUE;
--end HOLDX1;
--
--architecture behavioral of HOLDX1 is
--     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;
--
--     SIGNAL Y_ipd : std_ulogic := 'X';
--     SIGNAL io_wire : std_logic := 'X';
--     CONSTANT ResultMapping : VitalResultMapType := ('W', 'W', 'L', 'H');
--
--BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
-- functionality section
--        VITALBUF (io_wire, Y);
--        VITALBUF (Y, 
--                  io_wire,
--                  ( 0 ps, 0 ps),
--                  ResultMapping );
-- 
--end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX12 : entity is TRUE;
end INVX12;

architecture behavioral of INVX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX16 : entity is TRUE;
end INVX16;

architecture behavioral of INVX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX1 : entity is TRUE;
end INVX1;

architecture behavioral of INVX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX20 : entity is TRUE;
end INVX20;

architecture behavioral of INVX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX2 : entity is TRUE;
end INVX2;

architecture behavioral of INVX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX3 : entity is TRUE;
end INVX3;

architecture behavioral of INVX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX4 : entity is TRUE;
end INVX4;

architecture behavioral of INVX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVX8 : entity is TRUE;
end INVX8;

architecture behavioral of INVX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity INVXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of INVXL : entity is TRUE;
end INVXL;

architecture behavioral of INVXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
END BLOCK;

VITALBehavior : PROCESS (A_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINV(A_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFX1 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFX1 : entity is TRUE;
end JKFFX1;

architecture behavioral of JKFFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX1",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX1",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFX2 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFX2 : entity is TRUE;
end JKFFX2;

architecture behavioral of JKFFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX2",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX2",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFX4 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFX4 : entity is TRUE;
end JKFFX4;

architecture behavioral of JKFFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX4",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFX4",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFXL is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFXL : entity is TRUE;
end JKFFXL;

architecture behavioral of JKFFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFXL",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFXL",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFRX1 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFRX1 : entity is TRUE;
end JKFFRX1;

architecture behavioral of JKFFRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX1",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX1",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFRX2 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFRX2 : entity is TRUE;
end JKFFRX2;

architecture behavioral of JKFFRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX2",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX2",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFRX4 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFRX4 : entity is TRUE;
end JKFFRX4;

architecture behavioral of JKFFRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX4",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRX4",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFRXL is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFRXL : entity is TRUE;
end JKFFRXL;

architecture behavioral of JKFFRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRXL",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFRXL",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := '1';

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSX1 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSX1 : entity is TRUE;
end JKFFSX1;

architecture behavioral of JKFFSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX1",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX1",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSX2 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSX2 : entity is TRUE;
end JKFFSX2;

architecture behavioral of JKFFSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX2",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX2",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSX4 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSX4 : entity is TRUE;
end JKFFSX4;

architecture behavioral of JKFFSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX4",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSX4",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSXL is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSXL : entity is TRUE;
end JKFFSXL;

architecture behavioral of JKFFSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSXL",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSXL",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := '1';


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSRX1 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSRX1 : entity is TRUE;
end JKFFSRX1;

architecture behavioral of JKFFSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSRX2 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSRX2 : entity is TRUE;
end JKFFSRX2;

architecture behavioral of JKFFSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSRX4 is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSRX4 : entity is TRUE;
end JKFFSRX4;

architecture behavioral of JKFFSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: jkff.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity JKFFSRXL is

     generic ( tipd_J : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_K : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_J_CK : VitalDelayType := DefDummyIsd;
               tisd_K_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_J_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_J_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_J_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_J_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_K_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_K_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_K_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_K_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            J : in std_ulogic := 'U';
            K : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            CK : in std_ulogic := 'U');

     attribute VITAL_LEVEL0 of JKFFSRXL : entity is TRUE;
end JKFFSRXL;

architecture behavioral of JKFFSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL J_dly : std_ulogic := 'X';
     SIGNAL K_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL J_ipd : std_ulogic := 'X';
     SIGNAL K_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( J_ipd,  J, tipd_J );
          VitalWireDelay( K_ipd, K, tipd_K );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( J_dly, J_ipd, tisd_J_CK );
          VitalSignalDelay( K_dly, K_ipd, tisd_K_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (J_dly, K_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_J_CK : std_ulogic := '0';
     VARIABLE TimeMarker_J_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_K_CK : std_ulogic := '0';
     VARIABLE TimeMarker_K_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_jkff_n0 : std_logic_vector( 0 TO 5 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE S : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE xRN_dly : std_ulogic;

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SN_CK_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_CK_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_SN_CK,
                   Violation      => Tviol_SN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => J_dly,
                   TestSignalName => "J",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_J_CK_posedge_posedge,
                   SetupLow       => tsetup_J_CK_negedge_posedge,
                   HoldHigh       => thold_J_CK_negedge_posedge,
                   HoldLow        => thold_J_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_J_CK,
                   Violation      => Tviol_J_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => K_dly,
                   TestSignalName => "K",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_K_CK_posedge_posedge,
                   SetupLow       => tsetup_K_CK_negedge_posedge,
                   HoldHigh       => thold_K_CK_negedge_posedge,
                   HoldLow        => thold_K_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   TimingData     => TimeMarker_K_CK,
                   Violation      => Tviol_K_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/JKFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        Tviol_J_CK OR 
                        Tviol_K_CK OR 
                        PWviol_CK 
                      );

          xSN_dly := SN_dly;

          xRN_dly := RN_dly;


          VitalStateTable ( StateTable => udp_jkff,
                           DataIn => (NOTIFIER,J_dly,K_dly,CK_dly,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_jkff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          S := VitalBUF(xSN_dly );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             ( To_X01(S) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX2X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX2X1 : entity is TRUE;
end MX2X1;

architecture behavioral of MX2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX2X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX2X2 : entity is TRUE;
end MX2X2;

architecture behavioral of MX2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX2X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX2X4 : entity is TRUE;
end MX2X4;

architecture behavioral of MX2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX2XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX2XL : entity is TRUE;
end MX2XL;

architecture behavioral of MX2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX4X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX4X1 : entity is TRUE;
end MX4X1;

architecture behavioral of MX4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX4X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX4X2 : entity is TRUE;
end MX4X2;

architecture behavioral of MX4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX4X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX4X4 : entity is TRUE;
end MX4X4;

architecture behavioral of MX4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MX4XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MX4XL : entity is TRUE;
end MX4XL;

architecture behavioral of MX4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalBUF( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI2X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI2X1 : entity is TRUE;
end MXI2X1;

architecture behavioral of MXI2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI2X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI2X2 : entity is TRUE;
end MXI2X2;

architecture behavioral of MXI2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI2X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI2X4 : entity is TRUE;
end MXI2X4;

architecture behavioral of MXI2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI2XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
	       tpd_S0_Y_A_EQ_1_AN_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI2XL : entity is TRUE;
end MXI2XL;

architecture behavioral of MXI2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, S0_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux2( B_ipd, A_ipd,S0_ipd);
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1,
                             ((To_X01(A_ipd) /= '1') and (To_X01(B_ipd) /= '0'))),
                      3 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0,
                             ((To_X01(A_ipd) /= '0') and (To_X01(B_ipd) /= '1')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI4X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI4X1 : entity is TRUE;
end MXI4X1;

architecture behavioral of MXI4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI4X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI4X2 : entity is TRUE;
end MXI4X2;

architecture behavioral of MXI4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI4X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI4X4 : entity is TRUE;
end MXI4X4;

architecture behavioral of MXI4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: mux.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity MXI4XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_S1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
               );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U';
            S0 : in std_ulogic := 'U';
            S1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of MXI4XL : entity is TRUE;
end MXI4XL;

architecture behavioral of MXI4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL S0_ipd : std_ulogic := 'X';
     SIGNAL S1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( S0_ipd, S0, tipd_S0 );
          VitalWireDelay( S1_ipd, S1, tipd_S1 );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          n0 := VitalMux4((D_ipd & C_ipd & B_ipd & A_ipd),(S1_ipd  & S0_ipd));
     
          Y_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE ),
                      4 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_0_AN_B_EQ_1_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      5 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_A_EQ_1_AN_B_EQ_0_AN_S1_EQ_0,
                             ((To_X01(S1_ipd) /= '1') and (To_X01(B_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      6 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_0_AN_D_EQ_1_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(C_ipd) /= '1'))),
                      7 => ( S0_ipd'LAST_EVENT,
                             tpd_S0_Y_C_EQ_1_AN_D_EQ_0_AN_S1_EQ_1,
                             ((To_X01(S1_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(C_ipd) /= '0'))),
                      8 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_0_AN_C_EQ_1_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='0') and (To_X01(A_ipd) /= '1'))),
                      9 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_A_EQ_1_AN_C_EQ_0_AN_S0_EQ_0,
                             ((To_X01(S0_ipd) /= '1') and (To_X01(C_ipd) /='1') and (To_X01(A_ipd) /= '0'))),
                      10 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_0_AN_D_EQ_1_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='0') and (To_X01(B_ipd) /= '1'))),
                      11 => ( S1_ipd'LAST_EVENT,
                             tpd_S1_Y_B_EQ_1_AN_D_EQ_0_AN_S0_EQ_1,
                             ((To_X01(S0_ipd) /= '0') and (To_X01(D_ipd) /='1') and (To_X01(B_ipd) /= '0')))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2X1 : entity is TRUE;
end NAND2X1;

architecture behavioral of NAND2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2X2 : entity is TRUE;
end NAND2X2;

architecture behavioral of NAND2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2X4 : entity is TRUE;
end NAND2X4;

architecture behavioral of NAND2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2XL : entity is TRUE;
end NAND2XL;

architecture behavioral of NAND2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2BX1 : entity is TRUE;
end NAND2BX1;

architecture behavioral of NAND2BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2BX2 : entity is TRUE;
end NAND2BX2;

architecture behavioral of NAND2BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2BX4 : entity is TRUE;
end NAND2BX4;

architecture behavioral of NAND2BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND2BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND2BXL : entity is TRUE;
end NAND2BXL;

architecture behavioral of NAND2BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3X1 : entity is TRUE;
end NAND3X1;

architecture behavioral of NAND3X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3X2 : entity is TRUE;
end NAND3X2;

architecture behavioral of NAND3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3X4 : entity is TRUE;
end NAND3X4;

architecture behavioral of NAND3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3XL : entity is TRUE;
end NAND3XL;

architecture behavioral of NAND3XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3BX1 : entity is TRUE;
end NAND3BX1;

architecture behavioral of NAND3BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3BX2 : entity is TRUE;
end NAND3BX2;

architecture behavioral of NAND3BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3BX4 : entity is TRUE;
end NAND3BX4;

architecture behavioral of NAND3BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND3BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND3BXL : entity is TRUE;
end NAND3BXL;

architecture behavioral of NAND3BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4X1 : entity is TRUE;
end NAND4X1;

architecture behavioral of NAND4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4X2 : entity is TRUE;
end NAND4X2;

architecture behavioral of NAND4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4X4 : entity is TRUE;
end NAND4X4;

architecture behavioral of NAND4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4XL : entity is TRUE;
end NAND4XL;

architecture behavioral of NAND4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNAND4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BX1 : entity is TRUE;
end NAND4BX1;

architecture behavioral of NAND4BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BX2 : entity is TRUE;
end NAND4BX2;

architecture behavioral of NAND4BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BX4 : entity is TRUE;
end NAND4BX4;

architecture behavioral of NAND4BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BXL : entity is TRUE;
end NAND4BXL;

architecture behavioral of NAND4BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNAND4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BBX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BBX1 : entity is TRUE;
end NAND4BBX1;

architecture behavioral of NAND4BBX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNAND4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BBX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BBX2 : entity is TRUE;
end NAND4BBX2;

architecture behavioral of NAND4BBX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNAND4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BBX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BBX4 : entity is TRUE;
end NAND4BBX4;

architecture behavioral of NAND4BBX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNAND4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NAND4BBXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NAND4BBXL : entity is TRUE;
end NAND4BBXL;

architecture behavioral of NAND4BBXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNAND4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2X1 : entity is TRUE;
end NOR2X1;

architecture behavioral of NOR2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2X2 : entity is TRUE;
end NOR2X2;

architecture behavioral of NOR2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2X4 : entity is TRUE;
end NOR2X4;

architecture behavioral of NOR2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2XL : entity is TRUE;
end NOR2XL;

architecture behavioral of NOR2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2BX1 : entity is TRUE;
end NOR2BX1;

architecture behavioral of NOR2BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2BX2 : entity is TRUE;
end NOR2BX2;

architecture behavioral of NOR2BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2BX4 : entity is TRUE;
end NOR2BX4;

architecture behavioral of NOR2BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR2BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR2BXL : entity is TRUE;
end NOR2BXL;

architecture behavioral of NOR2BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR2(out1,B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3X1 : entity is TRUE;
end NOR3X1;

architecture behavioral of NOR3X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3X2 : entity is TRUE;
end NOR3X2;

architecture behavioral of NOR3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3X4 : entity is TRUE;
end NOR3X4;

architecture behavioral of NOR3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3XL : entity is TRUE;
end NOR3XL;

architecture behavioral of NOR3XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3BX1 : entity is TRUE;
end NOR3BX1;

architecture behavioral of NOR3BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3BX2 : entity is TRUE;
end NOR3BX2;

architecture behavioral of NOR3BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3BX4 : entity is TRUE;
end NOR3BX4;

architecture behavioral of NOR3BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR3BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR3BXL : entity is TRUE;
end NOR3BXL;

architecture behavioral of NOR3BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR3(out1,B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4X1 : entity is TRUE;
end NOR4X1;

architecture behavioral of NOR4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4X2 : entity is TRUE;
end NOR4X2;

architecture behavioral of NOR4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4X4 : entity is TRUE;
end NOR4X4;

architecture behavioral of NOR4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4XL : entity is TRUE;
end NOR4XL;

architecture behavioral of NOR4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalNOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BX1 : entity is TRUE;
end NOR4BX1;

architecture behavioral of NOR4BX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BX2 : entity is TRUE;
end NOR4BX2;

architecture behavioral of NOR4BX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BX4 : entity is TRUE;
end NOR4BX4;

architecture behavioral of NOR4BX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BXL : entity is TRUE;
end NOR4BXL;

architecture behavioral of NOR4BXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          Y_zd := VitalNOR4(out1,B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BBX1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BBX1 : entity is TRUE;
end NOR4BBX1;

architecture behavioral of NOR4BBX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNOR4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BBX2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BBX2 : entity is TRUE;
end NOR4BBX2;

architecture behavioral of NOR4BBX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNOR4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BBX4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BBX4 : entity is TRUE;
end NOR4BBX4;

architecture behavioral of NOR4BBX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNOR4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity NOR4BBXL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_AN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_AN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_BN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_BN_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            AN : in std_ulogic := 'U';
            BN : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of NOR4BBXL : entity is TRUE;
end NOR4BBXL;

architecture behavioral of NOR4BBXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL AN_ipd : std_ulogic := 'X';
     SIGNAL BN_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( AN_ipd, AN, tipd_AN );
          VitalWireDelay( BN_ipd, BN, tipd_BN );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (AN_ipd, BN_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE out1 : std_ulogic;
     VARIABLE out2 : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          out1 := VitalINV(AN_ipd);

          out2 := VitalINV(BN_ipd);

          Y_zd := VitalNOR4(out1,out2,C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( AN_ipd'LAST_EVENT,
                             tpd_AN_Y,
                             TRUE ),
                      1 => ( BN_ipd'LAST_EVENT,
                             tpd_BN_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI211X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI211X1 : entity is TRUE;
end OAI211X1;

architecture behavioral of OAI211X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI211X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI211X2 : entity is TRUE;
end OAI211X2;

architecture behavioral of OAI211X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI211X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI211X4 : entity is TRUE;
end OAI211X4;

architecture behavioral of OAI211X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI211XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI211XL : entity is TRUE;
end OAI211XL;

architecture behavioral of OAI211XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND3(outA, B0_ipd, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI21X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI21X1 : entity is TRUE;
end OAI21X1;

architecture behavioral of OAI21X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI21X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI21X2 : entity is TRUE;
end OAI21X2;

architecture behavioral of OAI21X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI21X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI21X4 : entity is TRUE;
end OAI21X4;

architecture behavioral of OAI21X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI21XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI21XL : entity is TRUE;
end OAI21XL;

architecture behavioral of OAI21XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI221X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI221X1 : entity is TRUE;
end OAI221X1;

architecture behavioral of OAI221X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI221X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI221X2 : entity is TRUE;
end OAI221X2;

architecture behavioral of OAI221X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI221X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI221X4 : entity is TRUE;
end OAI221X4;

architecture behavioral of OAI221X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI221XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI221XL : entity is TRUE;
end OAI221XL;

architecture behavioral of OAI221XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND3(outA, outB, C0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI222X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI222X1 : entity is TRUE;
end OAI222X1;

architecture behavioral of OAI222X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          outC := VitalOR2(C0_ipd, C1_ipd);

          Y_zd := VitalNAND3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI222X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI222X2 : entity is TRUE;
end OAI222X2;

architecture behavioral of OAI222X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          outC := VitalOR2(C0_ipd, C1_ipd);

          Y_zd := VitalNAND3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI222X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI222X4 : entity is TRUE;
end OAI222X4;

architecture behavioral of OAI222X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          outC := VitalOR2(C0_ipd, C1_ipd);

          Y_zd := VitalNAND3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI222XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            C0 : in std_ulogic := 'U';
            C1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI222XL : entity is TRUE;
end OAI222XL;

architecture behavioral of OAI222XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL C0_ipd : std_ulogic := 'X';
     SIGNAL C1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( C0_ipd, C0, tipd_C0 );
          VitalWireDelay( C1_ipd, C1, tipd_C1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd, C0_ipd, C1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          outC := VitalOR2(C0_ipd, C1_ipd);

          Y_zd := VitalNAND3(outA, outB, outC);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      4 => ( C0_ipd'LAST_EVENT,
                             tpd_C0_Y,
                             TRUE ),
                      5 => ( C1_ipd'LAST_EVENT,
                             tpd_C1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI22X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI22X1 : entity is TRUE;
end OAI22X1;

architecture behavioral of OAI22X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI22X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI22X2 : entity is TRUE;
end OAI22X2;

architecture behavioral of OAI22X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI22X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI22X4 : entity is TRUE;
end OAI22X4;

architecture behavioral of OAI22X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI22XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI22XL : entity is TRUE;
end OAI22XL;

architecture behavioral of OAI22XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR2(A0_ipd, A1_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB1X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB1X1 : entity is TRUE;
end OAI2BB1X1;

architecture behavioral of OAI2BB1X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB1X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB1X2 : entity is TRUE;
end OAI2BB1X2;

architecture behavioral of OAI2BB1X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB1X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB1X4 : entity is TRUE;
end OAI2BB1X4;

architecture behavioral of OAI2BB1X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB1XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB1XL : entity is TRUE;
end OAI2BB1XL;

architecture behavioral of OAI2BB1XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB2X1 : entity is TRUE;
end OAI2BB2X1;

architecture behavioral of OAI2BB2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB2X2 : entity is TRUE;
end OAI2BB2X2;

architecture behavioral of OAI2BB2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB2X4 : entity is TRUE;
end OAI2BB2X4;

architecture behavioral of OAI2BB2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI2BB2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1N : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1N_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0N : in std_ulogic := 'U';
            A1N : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI2BB2XL : entity is TRUE;
end OAI2BB2XL;

architecture behavioral of OAI2BB2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0N_ipd : std_ulogic := 'X';
     SIGNAL A1N_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0N_ipd, A0N, tipd_A0N );
          VitalWireDelay( A1N_ipd, A1N, tipd_A1N );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0N_ipd, A1N_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;
     VARIABLE A0X_ipd   : std_ulogic;
     VARIABLE A1X_ipd   : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          A0X_ipd := VitalINV(A0N_ipd);

          A1X_ipd := VitalINV(A1N_ipd);

          outA := VitalOR2(A0X_ipd, A1X_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0N_ipd'LAST_EVENT,
                             tpd_A0N_Y,
                             TRUE ),
                      1 => ( A1N_ipd'LAST_EVENT,
                             tpd_A1N_Y,
                             TRUE ),
                      2 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      3 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI31X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI31X1 : entity is TRUE;
end OAI31X1;

architecture behavioral of OAI31X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI31X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI31X2 : entity is TRUE;
end OAI31X2;

architecture behavioral of OAI31X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI31X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI31X4 : entity is TRUE;
end OAI31X4;

architecture behavioral of OAI31X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI31XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI31XL : entity is TRUE;
end OAI31XL;

architecture behavioral of OAI31XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          Y_zd := VitalNAND2(outA, B0_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI32X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI32X1 : entity is TRUE;
end OAI32X1;

architecture behavioral of OAI32X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI32X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI32X2 : entity is TRUE;
end OAI32X2;

architecture behavioral of OAI32X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI32X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI32X4 : entity is TRUE;
end OAI32X4;

architecture behavioral of OAI32X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI32XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI32XL : entity is TRUE;
end OAI32XL;

architecture behavioral of OAI32XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR2(B0_ipd, B1_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI33X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI33X1 : entity is TRUE;
end OAI33X1;

architecture behavioral of OAI33X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI33X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI33X2 : entity is TRUE;
end OAI33X2;

architecture behavioral of OAI33X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI33X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI33X4 : entity is TRUE;
end OAI33X4;

architecture behavioral of OAI33X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: aoi.genpp,v 1.6 2002/01/28 22:03:18 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OAI33XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_A2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B0 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B0_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B1 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B1_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B2 : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B2_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A0 : in std_ulogic := 'U';
            A1 : in std_ulogic := 'U';
            A2 : in std_ulogic := 'U';
            B0 : in std_ulogic := 'U';
            B1 : in std_ulogic := 'U';
            B2 : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OAI33XL : entity is TRUE;
end OAI33XL;

architecture behavioral of OAI33XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A0_ipd : std_ulogic := 'X';
     SIGNAL A1_ipd : std_ulogic := 'X';
     SIGNAL A2_ipd : std_ulogic := 'X';
     SIGNAL B0_ipd : std_ulogic := 'X';
     SIGNAL B1_ipd : std_ulogic := 'X';
     SIGNAL B2_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A0_ipd, A0, tipd_A0 );
          VitalWireDelay( A1_ipd, A1, tipd_A1 );
          VitalWireDelay( A2_ipd, A2, tipd_A2 );
          VitalWireDelay( B0_ipd, B0, tipd_B0 );
          VitalWireDelay( B1_ipd, B1, tipd_B1 );
          VitalWireDelay( B2_ipd, B2, tipd_B2 );
END BLOCK;

VITALBehavior : PROCESS (A0_ipd, A1_ipd, A2_ipd, B0_ipd, B1_ipd, B2_ipd)


     -- functionality section variables
     VARIABLE outA : std_ulogic;
     VARIABLE outB : std_ulogic;
     VARIABLE outC : std_ulogic;
     VARIABLE outD : std_ulogic;
     VARIABLE outA1 : std_ulogic;
     VARIABLE outB1 : std_ulogic;
     VARIABLE outC1 : std_ulogic;
     VARIABLE outD1 : std_ulogic;
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          outA := VitalOR3(A0_ipd, A1_ipd, A2_ipd);

          outB := VitalOR3(B0_ipd, B1_ipd, B2_ipd);

          Y_zd := VitalNAND2(outA, outB);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A0_ipd'LAST_EVENT,
                             tpd_A0_Y,
                             TRUE ),
                      1 => ( A1_ipd'LAST_EVENT,
                             tpd_A1_Y,
                             TRUE ),
                      2 => ( A2_ipd'LAST_EVENT,
                             tpd_A2_Y,
                             TRUE ),
                      3 => ( B0_ipd'LAST_EVENT,
                             tpd_B0_Y,
                             TRUE ),
                      4 => ( B1_ipd'LAST_EVENT,
                             tpd_B1_Y,
                             TRUE ),
                      5 => ( B2_ipd'LAST_EVENT,
                             tpd_B2_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR2X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR2X1 : entity is TRUE;
end OR2X1;

architecture behavioral of OR2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR2X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR2X2 : entity is TRUE;
end OR2X2;

architecture behavioral of OR2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR2X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR2X4 : entity is TRUE;
end OR2X4;

architecture behavioral of OR2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR2XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR2XL : entity is TRUE;
end OR2XL;

architecture behavioral of OR2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR2(A_ipd, B_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR3X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR3X1 : entity is TRUE;
end OR3X1;

architecture behavioral of OR3X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR3X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR3X2 : entity is TRUE;
end OR3X2;

architecture behavioral of OR3X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR3X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR3X4 : entity is TRUE;
end OR3X4;

architecture behavioral of OR3X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR3XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR3XL : entity is TRUE;
end OR3XL;

architecture behavioral of OR3XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR3(A_ipd, B_ipd, C_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR4X1 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR4X1 : entity is TRUE;
end OR4X1;

architecture behavioral of OR4X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR4X2 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR4X2 : entity is TRUE;
end OR4X2;

architecture behavioral of OR4X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR4X4 is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR4X4 : entity is TRUE;
end OR4X4;

architecture behavioral of OR4X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: comb.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity OR4XL is

     generic ( 
               XOn          : BOOLEAN := DefCombSpikeXOn;
               MsgOn        : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING  := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_C : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_C_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_D_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
             );

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U';
            C : in std_ulogic := 'U';
            D : in std_ulogic := 'U'
          );

     attribute VITAL_LEVEL0 of OR4XL : entity is TRUE;
end OR4XL;

architecture behavioral of OR4XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';
     SIGNAL C_ipd : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
          VitalWireDelay( C_ipd, C, tipd_C );
          VitalWireDelay( D_ipd, D, tipd_D );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd, C_ipd, D_ipd)

     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n1 : std_ulogic;
    

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalOR4(A_ipd, B_ipd, C_ipd, D_ipd);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y,
                             TRUE ),
                      1 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y,
                             TRUE ),
                      2 => ( C_ipd'LAST_EVENT,
                             tpd_C_Y,
                             TRUE ),
                      3 => ( D_ipd'LAST_EVENT,
                             tpd_D_Y,
                             TRUE )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATX1 is

     generic ( 
               tipd_R : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_R_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_R_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_R_posedge : VitalDelayType := DefDummyWidth;
               tipd_S : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_S_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_S_posedge : VitalDelayType := DefDummyWidth;
               thold_R_S_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               thold_S_R_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            R : in std_ulogic := 'U';
            S : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATX1 : entity is TRUE;
end RSLATX1;

architecture behavioral of RSLATX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL R_ipd : std_ulogic := 'X';
     SIGNAL S_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( R_ipd, R, tipd_R );
          VitalWireDelay( S_ipd, S, tipd_S );
     END BLOCK;


     VITALBehavior : PROCESS (R_ipd, S_ipd)

          -- timing check section variables
          VARIABLE Tviol_S_R_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_S_R_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_R_S_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_R_S_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_S_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_S_posedge : VitalPeriodDataType;
          VARIABLE PWviol_R_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_R_posedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslat_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslat_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   RefSignal      => S_ipd,
                   RefSignalName  => "S",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_S_R_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX1",
                   TimingData     => TimeMarker_S_R_negedge,
                   Violation      => Tviol_S_R_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   RefSignal      => R_ipd,
                   RefSignalName  => "R",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_R_S_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX1",
                   TimingData     => TimeMarker_R_S_negedge,
                   Violation      => Tviol_R_S_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_S_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_S_posedge,
                   Violation      => PWviol_S_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_R_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_R_posedge,
                   Violation      => PWviol_R_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_S_R_negedge OR Tviol_R_S_negedge OR PWviol_S_posedge OR PWviol_R_posedge );

     VitalStateTable ( StateTable => udp_rslat_out,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslat_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslat_out_n,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslat_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_Q,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_QN,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATX2 is

     generic ( 
               tipd_R : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_R_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_R_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_R_posedge : VitalDelayType := DefDummyWidth;
               tipd_S : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_S_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_S_posedge : VitalDelayType := DefDummyWidth;
               thold_R_S_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               thold_S_R_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            R : in std_ulogic := 'U';
            S : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATX2 : entity is TRUE;
end RSLATX2;

architecture behavioral of RSLATX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL R_ipd : std_ulogic := 'X';
     SIGNAL S_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( R_ipd, R, tipd_R );
          VitalWireDelay( S_ipd, S, tipd_S );
     END BLOCK;


     VITALBehavior : PROCESS (R_ipd, S_ipd)

          -- timing check section variables
          VARIABLE Tviol_S_R_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_S_R_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_R_S_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_R_S_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_S_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_S_posedge : VitalPeriodDataType;
          VARIABLE PWviol_R_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_R_posedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslat_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslat_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   RefSignal      => S_ipd,
                   RefSignalName  => "S",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_S_R_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX2",
                   TimingData     => TimeMarker_S_R_negedge,
                   Violation      => Tviol_S_R_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   RefSignal      => R_ipd,
                   RefSignalName  => "R",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_R_S_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX2",
                   TimingData     => TimeMarker_R_S_negedge,
                   Violation      => Tviol_R_S_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_S_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_S_posedge,
                   Violation      => PWviol_S_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_R_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_R_posedge,
                   Violation      => PWviol_R_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_S_R_negedge OR Tviol_R_S_negedge OR PWviol_S_posedge OR PWviol_R_posedge );

     VitalStateTable ( StateTable => udp_rslat_out,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslat_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslat_out_n,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslat_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_Q,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_QN,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATX4 is

     generic ( 
               tipd_R : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_R_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_R_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_R_posedge : VitalDelayType := DefDummyWidth;
               tipd_S : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_S_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_S_posedge : VitalDelayType := DefDummyWidth;
               thold_R_S_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               thold_S_R_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            R : in std_ulogic := 'U';
            S : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATX4 : entity is TRUE;
end RSLATX4;

architecture behavioral of RSLATX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL R_ipd : std_ulogic := 'X';
     SIGNAL S_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( R_ipd, R, tipd_R );
          VitalWireDelay( S_ipd, S, tipd_S );
     END BLOCK;


     VITALBehavior : PROCESS (R_ipd, S_ipd)

          -- timing check section variables
          VARIABLE Tviol_S_R_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_S_R_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_R_S_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_R_S_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_S_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_S_posedge : VitalPeriodDataType;
          VARIABLE PWviol_R_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_R_posedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslat_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslat_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   RefSignal      => S_ipd,
                   RefSignalName  => "S",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_S_R_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX4",
                   TimingData     => TimeMarker_S_R_negedge,
                   Violation      => Tviol_S_R_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   RefSignal      => R_ipd,
                   RefSignalName  => "R",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_R_S_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATX4",
                   TimingData     => TimeMarker_R_S_negedge,
                   Violation      => Tviol_R_S_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_S_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_S_posedge,
                   Violation      => PWviol_S_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_R_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_R_posedge,
                   Violation      => PWviol_R_posedge,
                   HeaderMsg      => InstancePath & "/RSLATX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_S_R_negedge OR Tviol_R_S_negedge OR PWviol_S_posedge OR PWviol_R_posedge );

     VitalStateTable ( StateTable => udp_rslat_out,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslat_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslat_out_n,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslat_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_Q,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_QN,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATXL is

     generic ( 
               tipd_R : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_R_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_R_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_R_posedge : VitalDelayType := DefDummyWidth;
               tipd_S : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_S_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_S_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_S_posedge : VitalDelayType := DefDummyWidth;
               thold_R_S_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               thold_S_R_negedge_negedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            R : in std_ulogic := 'U';
            S : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATXL : entity is TRUE;
end RSLATXL;

architecture behavioral of RSLATXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL R_ipd : std_ulogic := 'X';
     SIGNAL S_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( R_ipd, R, tipd_R );
          VitalWireDelay( S_ipd, S, tipd_S );
     END BLOCK;


     VITALBehavior : PROCESS (R_ipd, S_ipd)

          -- timing check section variables
          VARIABLE Tviol_S_R_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_S_R_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_R_S_negedge : std_ulogic := '0';
          VARIABLE TimeMarker_R_S_negedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_S_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_S_posedge : VitalPeriodDataType;
          VARIABLE PWviol_R_posedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_R_posedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslat_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslat_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   RefSignal      => S_ipd,
                   RefSignalName  => "S",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_S_R_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATXL",
                   TimingData     => TimeMarker_S_R_negedge,
                   Violation      => Tviol_S_R_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   RefSignal      => R_ipd,
                   RefSignalName  => "R",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => thold_R_S_negedge_negedge,
                   HoldLow        => 0 ps,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/RSLATXL",
                   TimingData     => TimeMarker_R_S_negedge,
                   Violation      => Tviol_R_S_negedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => S_ipd,
                   TestSignalName => "S",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_S_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_S_posedge,
                   Violation      => PWviol_S_posedge,
                   HeaderMsg      => InstancePath & "/RSLATXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => R_ipd,
                   TestSignalName => "R",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_R_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_R_posedge,
                   Violation      => PWviol_R_posedge,
                   HeaderMsg      => InstancePath & "/RSLATXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_S_R_negedge OR Tviol_R_S_negedge OR PWviol_S_posedge OR PWviol_R_posedge );

     VitalStateTable ( StateTable => udp_rslat_out,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslat_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslat_out_n,
                        DataIn => (NOTIFIER, R_ipd, S_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslat_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_Q,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( R_ipd'LAST_EVENT,
                             tpd_R_QN,
                             TRUE ),
                      1 => ( S_ipd'LAST_EVENT,
                             tpd_S_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATNX1 is

     generic ( 
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            RN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATNX1 : entity is TRUE;
end RSLATNX1;

architecture behavioral of RSLATNX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( RN_ipd, RN, tipd_RN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
     END BLOCK;


     VITALBehavior : PROCESS (RN_ipd, SN_ipd)

          -- timing check section variables
          VARIABLE Tviol_SN_RN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_SN_RN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_RN_SN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_RN_SN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_SN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
          VARIABLE PWviol_RN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslatn_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslatn_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   RefSignal      => SN_ipd,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX1",
                   TimingData     => TimeMarker_SN_RN_posedge,
                   Violation      => Tviol_SN_RN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   RefSignal      => RN_ipd,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX1",
                   TimingData     => TimeMarker_RN_SN_posedge,
                   Violation      => Tviol_RN_SN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_SN_RN_posedge OR Tviol_RN_SN_posedge OR PWviol_SN_negedge OR PWviol_RN_negedge );

     VitalStateTable ( StateTable => udp_rslatn_out,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslatn_out_n,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATNX2 is

     generic ( 
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            RN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATNX2 : entity is TRUE;
end RSLATNX2;

architecture behavioral of RSLATNX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( RN_ipd, RN, tipd_RN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
     END BLOCK;


     VITALBehavior : PROCESS (RN_ipd, SN_ipd)

          -- timing check section variables
          VARIABLE Tviol_SN_RN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_SN_RN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_RN_SN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_RN_SN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_SN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
          VARIABLE PWviol_RN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslatn_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslatn_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   RefSignal      => SN_ipd,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX2",
                   TimingData     => TimeMarker_SN_RN_posedge,
                   Violation      => Tviol_SN_RN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   RefSignal      => RN_ipd,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX2",
                   TimingData     => TimeMarker_RN_SN_posedge,
                   Violation      => Tviol_RN_SN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_SN_RN_posedge OR Tviol_RN_SN_posedge OR PWviol_SN_negedge OR PWviol_RN_negedge );

     VitalStateTable ( StateTable => udp_rslatn_out,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslatn_out_n,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATNX4 is

     generic ( 
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            RN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATNX4 : entity is TRUE;
end RSLATNX4;

architecture behavioral of RSLATNX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( RN_ipd, RN, tipd_RN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
     END BLOCK;


     VITALBehavior : PROCESS (RN_ipd, SN_ipd)

          -- timing check section variables
          VARIABLE Tviol_SN_RN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_SN_RN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_RN_SN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_RN_SN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_SN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
          VARIABLE PWviol_RN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslatn_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslatn_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   RefSignal      => SN_ipd,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX4",
                   TimingData     => TimeMarker_SN_RN_posedge,
                   Violation      => Tviol_SN_RN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   RefSignal      => RN_ipd,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNX4",
                   TimingData     => TimeMarker_RN_SN_posedge,
                   Violation      => Tviol_RN_SN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_SN_RN_posedge OR Tviol_RN_SN_posedge OR PWviol_SN_negedge OR PWviol_RN_negedge );

     VitalStateTable ( StateTable => udp_rslatn_out,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslatn_out_n,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: rslat.genpp,v 1.3 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity RSLATNXL is

     generic ( 
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            RN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q  : out std_ulogic;
            QN : out std_ulogic
          );

     attribute VITAL_LEVEL0 of RSLATNXL : entity is TRUE;
end RSLATNXL;

architecture behavioral of RSLATNXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL RN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

     ---------------------------------------------------
     -- Input Path Delays
     ---------------------------------------------------
     WIREDELAY : BLOCK
     BEGIN
          VitalWireDelay( RN_ipd, RN, tipd_RN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
     END BLOCK;


     VITALBehavior : PROCESS (RN_ipd, SN_ipd)

          -- timing check section variables
          VARIABLE Tviol_SN_RN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_SN_RN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE Tviol_RN_SN_posedge : std_ulogic := '0';
          VARIABLE TimeMarker_RN_SN_posedge : VitalTimingDataType := VitalTimingDataInit;
          VARIABLE PWviol_SN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
          VARIABLE PWviol_RN_negedge : std_ulogic := '0';
          VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;

          -- functionality section variables
          VARIABLE qint : std_ulogic;
          VARIABLE qint_vec : std_logic_vector( 1 TO 1 );
          VARIABLE qund : std_ulogic;
          VARIABLE qund_vec : std_logic_vector( 1 TO 1 );
          VARIABLE QN_zd : std_ulogic;
          VARIABLE Q_zd : std_ulogic;
          VARIABLE NOTIFIER : std_ulogic := '0';
          VARIABLE PrevData_udp_rslatn_out: std_logic_vector( 0 TO 2 );
          VARIABLE PrevData_udp_rslatn_out_n: std_logic_vector( 0 TO 2 );

          -- path delay section variables
          VARIABLE Q_GlitchData : VitalGlitchDataType;
          VARIABLE QN_GlitchData : VitalGlitchDataType;

     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   RefSignal      => SN_ipd,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNXL",
                   TimingData     => TimeMarker_SN_RN_posedge,
                   Violation      => Tviol_SN_RN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   RefSignal      => RN_ipd,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/RSLATNXL",
                   TimingData     => TimeMarker_RN_SN_posedge,
                   Violation      => Tviol_RN_SN_posedge,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_ipd,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_ipd,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/RSLATNXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


-- functionality section
          NOTIFIER := ( Tviol_SN_RN_posedge OR Tviol_RN_SN_posedge OR PWviol_SN_negedge OR PWviol_RN_negedge );

     VitalStateTable ( StateTable => udp_rslatn_out,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qint_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out );
     qint := qint_vec(1);

     Q_zd := VitalBUF( qint );

     VitalStateTable ( StateTable => udp_rslatn_out_n,
                        DataIn => (NOTIFIER, RN_ipd, SN_ipd),
                        NumStates => 1,
                           Result => qund_vec,
                   PreviousDataIn => PrevData_udp_rslatn_out_n );
     qund := qund_vec(1);

     QN_zd := VitalBUF( qund );


          ---------------------------------------------------
          -- Path Delay section
          ---------------------------------------------------

          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( RN_ipd'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE ),
                      1 => ( SN_ipd'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);


     END PROCESS;

end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFX1 : entity is TRUE;
end SDFFX1;

architecture behavioral of SDFFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFX2 : entity is TRUE;
end SDFFX2;

architecture behavioral of SDFFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFX4 : entity is TRUE;
end SDFFX4;

architecture behavioral of SDFFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFXL : entity is TRUE;
end SDFFXL;

architecture behavioral of SDFFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFHQX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFHQX1 : entity is TRUE;
end SDFFHQX1;

architecture behavioral of SDFFHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFHQX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFHQX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFHQX2 : entity is TRUE;
end SDFFHQX2;

architecture behavioral of SDFFHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFHQX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFHQX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFHQX4 : entity is TRUE;
end SDFFHQX4;

architecture behavioral of SDFFHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFHQX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFHQXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFHQXL : entity is TRUE;
end SDFFHQXL;

architecture behavioral of SDFFHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFHQXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFHQXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNX1 : entity is TRUE;
end SDFFNX1;

architecture behavioral of SDFFNX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX1",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX1",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNX2 : entity is TRUE;
end SDFFNX2;

architecture behavioral of SDFFNX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX2",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX2",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNX4 : entity is TRUE;
end SDFFNX4;

architecture behavioral of SDFFNX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX4",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNX4",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNXL : entity is TRUE;
end SDFFNXL;

architecture behavioral of SDFFNXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNXL",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNXL",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNRX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNRX1 : entity is TRUE;
end SDFFNRX1;

architecture behavioral of SDFFNRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNRX1",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX1",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX1",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNRX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNRX2 : entity is TRUE;
end SDFFNRX2;

architecture behavioral of SDFFNRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNRX2",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX2",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX2",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNRX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNRX4 : entity is TRUE;
end SDFFNRX4;

architecture behavioral of SDFFNRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNRX4",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX4",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRX4",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNRXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNRXL : entity is TRUE;
end SDFFNRXL;

architecture behavioral of SDFFNRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNRXL",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRXL",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNRXL",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSX1 : entity is TRUE;
end SDFFNSX1;

architecture behavioral of SDFFNSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSX1",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX1",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX1",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSX2 : entity is TRUE;
end SDFFNSX2;

architecture behavioral of SDFFNSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSX2",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX2",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX2",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSX4 : entity is TRUE;
end SDFFNSX4;

architecture behavioral of SDFFNSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSX4",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX4",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSX4",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSXL : entity is TRUE;
end SDFFNSXL;

architecture behavioral of SDFFNSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSXL",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSXL",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSXL",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSRX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSRX1 : entity is TRUE;
end SDFFNSRX1;

architecture behavioral of SDFFNSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX1",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX1",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSRX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSRX2 : entity is TRUE;
end SDFFNSRX2;

architecture behavioral of SDFFNSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX2",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX2",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSRX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSRX4 : entity is TRUE;
end SDFFNSRX4;

architecture behavioral of SDFFNSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX4",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRX4",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFNSRXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CKN : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CKN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CKN : VitalDelayType := DefDummyIsd;
               tisd_SE_CKN : VitalDelayType := DefDummyIsd;
               ticd_CKN : VitalDelayType := DefDummyIcd;
               tpd_CKN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SI_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SI_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CKN_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_SE_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_SE_CKN_negedge_negedge : VitalDelayType := DefDummyHold;
               tpw_CKN_negedge : VitalDelayType := DefDummyWidth;
               tpw_CKN_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CKN : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CKN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CKN_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_CKN_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CKN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CKN : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFNSRXL : entity is TRUE;
end SDFFNSRXL;

architecture behavioral of SDFFNSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CKN_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CKN_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CKN_ipd, CKN, tipd_CKN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CKN );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CKN );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CKN );
          VitalSignalDelay( CKN_dly, CKN_ipd, ticd_CKN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CKN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CKN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CKN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_D_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CKN : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CKN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CKN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CKN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_RN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRXL",
                    TimingData     => TimeMarker_RN_CKN,
                    Violation      => Tviol_RN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CKN_dly,
                    RefSignalName  => "CKN",
                    SetupHigh      => tsetup_SN_CKN_posedge_negedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CKN_posedge_negedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'F',
                    HeaderMsg      => InstancePath & "/SDFFNSRXL",
                    TimingData     => TimeMarker_SN_CKN,
                    Violation      => Tviol_SN_CKN,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_D_CKN_posedge_negedge,
                   SetupLow       => tsetup_D_CKN_negedge_negedge,
                   HoldHigh       => thold_D_CKN_negedge_negedge,
                   HoldLow        => thold_D_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   TimingData     => TimeMarker_D_CKN,
                   Violation      => Tviol_D_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SI_CKN_posedge_negedge,
                   SetupLow       => tsetup_SI_CKN_negedge_negedge,
                   HoldHigh       => thold_SI_CKN_negedge_negedge,
                   HoldLow        => thold_SI_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   TimingData     => TimeMarker_SI_CKN,
                   Violation      => Tviol_SI_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CKN_dly,
                   RefSignalName  => "CKN",
                   SetupHigh      => tsetup_SE_CKN_posedge_negedge,
                   SetupLow       => tsetup_SE_CKN_negedge_negedge,
                   HoldHigh       => thold_SE_CKN_negedge_negedge,
                   HoldLow        => thold_SE_CKN_posedge_negedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   TimingData     => TimeMarker_SE_CKN,
                   Violation      => Tviol_SE_CKN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CKN_dly,
                   TestSignalName => "CKN",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CKN_posedge,
                   PulseWidthLow  => tpw_CKN_negedge,
                   PeriodData     => PeriodCheckInfo_CKN,
                   Violation      => PWviol_CKN,
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CKN OR 
                        Tviol_SI_CKN OR 
                        Tviol_SE_CKN OR 
                        Tviol_SN_CKN OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CKN OR 
                        PWviol_RN_negedge OR
                        PWviol_CKN  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalINV(CKN_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CKN_dly'LAST_EVENT,
                             tpd_CKN_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRX1 : entity is TRUE;
end SDFFRX1;

architecture behavioral of SDFFRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRX1",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRX2 : entity is TRUE;
end SDFFRX2;

architecture behavioral of SDFFRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRX2",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRX4 : entity is TRUE;
end SDFFRX4;

architecture behavioral of SDFFRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRX4",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRXL : entity is TRUE;
end SDFFRXL;

architecture behavioral of SDFFRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRXL",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRHQX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRHQX1 : entity is TRUE;
end SDFFRHQX1;

architecture behavioral of SDFFRHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRHQX1",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRHQX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRHQX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRHQX2 : entity is TRUE;
end SDFFRHQX2;

architecture behavioral of SDFFRHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRHQX2",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRHQX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRHQX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRHQX4 : entity is TRUE;
end SDFFRHQX4;

architecture behavioral of SDFFRHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRHQX4",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRHQX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFRHQXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFRHQXL : entity is TRUE;
end SDFFRHQXL;

architecture behavioral of SDFFRHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFRHQXL",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFRHQXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFRHQXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSX1 : entity is TRUE;
end SDFFSX1;

architecture behavioral of SDFFSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSX1",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSX2 : entity is TRUE;
end SDFFSX2;

architecture behavioral of SDFFSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSX2",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSX4 : entity is TRUE;
end SDFFSX4;

architecture behavioral of SDFFSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSX4",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSXL : entity is TRUE;
end SDFFSXL;

architecture behavioral of SDFFSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSXL",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSHQX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSHQX1 : entity is TRUE;
end SDFFSHQX1;

architecture behavioral of SDFFSHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSHQX1",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSHQX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSHQX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSHQX2 : entity is TRUE;
end SDFFSHQX2;

architecture behavioral of SDFFSHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSHQX2",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSHQX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSHQX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSHQX4 : entity is TRUE;
end SDFFSHQX4;

architecture behavioral of SDFFSHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSHQX4",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSHQX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSHQXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSHQXL : entity is TRUE;
end SDFFSHQXL;

architecture behavioral of SDFFSHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSHQXL",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSHQXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSHQXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := '1';

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRX1 : entity is TRUE;
end SDFFSRX1;

architecture behavioral of SDFFSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX1",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX1",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRX2 : entity is TRUE;
end SDFFSRX2;

architecture behavioral of SDFFSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX2",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX2",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRX4 : entity is TRUE;
end SDFFSRX4;

architecture behavioral of SDFFSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX4",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRX4",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRXL : entity is TRUE;
end SDFFSRXL;

architecture behavioral of SDFFSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRXL",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRXL",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRHQX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRHQX1 : entity is TRUE;
end SDFFSRHQX1;

architecture behavioral of SDFFSRHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRHQX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRHQX2 : entity is TRUE;
end SDFFSRHQX2;

architecture behavioral of SDFFSRHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRHQX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRHQX4 : entity is TRUE;
end SDFFSRHQX4;

architecture behavioral of SDFFSRHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFSRHQXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tisd_SN_CK : VitalDelayType := DefDummyIsd;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_SN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFSRHQXL : entity is TRUE;
end SDFFSRHQXL;

architecture behavioral of SDFFSRHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );


                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

                VitalSetupHoldCheck (
                    TestSignal     => SN_dly,
                    TestSignalName => "SN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_SN_CK_posedge_posedge,
                    SetupLow       => 0 ps,
                    HoldHigh       => 0 ps,
                    HoldLow        => thold_SN_CK_posedge_posedge,
                    CheckEnabled   => TRUE,
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                    TimingData     => TimeMarker_SN_CK,
                    Violation      => Tviol_SN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/SDFFSRHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_SN_CK OR 
                        PWviol_SN_negedge OR 
                        Tviol_RN_CK OR 
                        PWviol_RN_negedge OR
                        PWviol_CK  
                       );

          SNx_dly := SN_dly;

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          n1 := VitalTruthTable ( TruthTable => udp_mux,
                                  DataIn => (D_dly,SI_dly,SE_dly) );

          VitalStateTable ( StateTable => udp_dff,
                           DataIn => (NOTIFIER,n1,intclk,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_dff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             To_X01(SandR) /= '0' 
                           ),
                      1 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFTRX1 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFTRX1 : entity is TRUE;
end SDFFTRX1;

architecture behavioral of SDFFTRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE RNcheck : std_ulogic;
     VARIABLE E_dly : std_ulogic;
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => tsetup_RN_CK_negedge_posedge,
                    HoldHigh       => thold_RN_CK_negedge_posedge,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => To_X01(RNcheck) /= '0',
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFTRX1",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFTRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          E_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);
 
          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          RNcheck := VitalBUF(SNx_dly);
 
          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFTRX2 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFTRX2 : entity is TRUE;
end SDFFTRX2;

architecture behavioral of SDFFTRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE RNcheck : std_ulogic;
     VARIABLE E_dly : std_ulogic;
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => tsetup_RN_CK_negedge_posedge,
                    HoldHigh       => thold_RN_CK_negedge_posedge,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => To_X01(RNcheck) /= '0',
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFTRX2",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFTRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          E_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);
 
          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          RNcheck := VitalBUF(SNx_dly);
 
          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFTRX4 is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFTRX4 : entity is TRUE;
end SDFFTRX4;

architecture behavioral of SDFFTRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE RNcheck : std_ulogic;
     VARIABLE E_dly : std_ulogic;
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => tsetup_RN_CK_negedge_posedge,
                    HoldHigh       => thold_RN_CK_negedge_posedge,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => To_X01(RNcheck) /= '0',
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFTRX4",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFTRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          E_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);
 
          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          RNcheck := VitalBUF(SNx_dly);
 
          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: sdff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SDFFTRXL is

     generic (
               tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);

               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( 
            D : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            QN : out std_ulogic;
            Q : out std_ulogic
          );

     attribute VITAL_LEVEL0 of SDFFTRXL : entity is TRUE;
end SDFFTRXL;

architecture behavioral of SDFFTRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_dff_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE intclk : std_ulogic;
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE RNcheck : std_ulogic;
     VARIABLE E_dly : std_ulogic;
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandSE : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE SandRandSEb : std_ulogic;
     VARIABLE DxorSD : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

                VitalSetupHoldCheck (
                    TestSignal     => RN_dly,
                    TestSignalName => "RN",
                    RefSignal      => CK_dly,
                    RefSignalName  => "CK",
                    SetupHigh      => tsetup_RN_CK_posedge_posedge,
                    SetupLow       => tsetup_RN_CK_negedge_posedge,
                    HoldHigh       => thold_RN_CK_negedge_posedge,
                    HoldLow        => thold_RN_CK_posedge_posedge,
                    CheckEnabled   => To_X01(RNcheck) /= '0',
                    RefTransition  => 'R',
                    HeaderMsg      => InstancePath & "/SDFFTRXL",
                    TimingData     => TimeMarker_RN_CK,
                    Violation      => Tviol_RN_CK,
                    XOn            => DefSeqXOn,
                    MsgOn          => DefSeqMsgOn,
                    MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSEb) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(SandRandSE) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SDFFTRXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SDFFTRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                        Tviol_D_CK OR 
                        Tviol_SI_CK OR 
                        Tviol_SE_CK OR 
                        Tviol_RN_CK OR 
                        PWviol_CK  
                       );

          SNx_dly := '1';

          RNx_dly := RN_dly;

          intclk := VitalBUF(CK_dly);

          E_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);
 
          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandSE := VitalAND2(SandR,SE_dly);

          SEb := VitalINV( SE_dly );

          SandRandSEb := VitalAND2(SandR,SEb);

          DxorSD := VitalXOR2(D_dly,SI_dly);

          flag := VitalAND2(DxorSD,SandR);

          RNcheck := VitalBUF(SNx_dly);
 
          QN_zd := VitalINV( n0 );


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFHQX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFHQX1 : entity is TRUE;
end SEDFFHQX1;

architecture behavioral of SEDFFHQX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX1",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFHQX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFHQX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFHQX2 : entity is TRUE;
end SEDFFHQX2;

architecture behavioral of SEDFFHQX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX2",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFHQX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFHQX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFHQX4 : entity is TRUE;
end SEDFFHQX4;

architecture behavioral of SEDFFHQX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX4",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFHQX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFHQXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFHQXL : entity is TRUE;
end SEDFFHQXL;

architecture behavioral of SEDFFHQXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQXL",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFHQXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFHQXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFX1 : entity is TRUE;
end SEDFFX1;

architecture behavioral of SEDFFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX1",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFX2 : entity is TRUE;
end SEDFFX2;

architecture behavioral of SEDFFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX2",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFX4 : entity is TRUE;
end SEDFFX4;

architecture behavioral of SEDFFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX4",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFXL : entity is TRUE;
end SEDFFXL;

architecture behavioral of SEDFFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedff_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFXL",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := '1';

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedff,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedff_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          NoSetReset := VitalAND2(RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             ( To_X01(NoSetReset) ) /= '0' 
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFTRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFTRX1 : entity is TRUE;
end SEDFFTRX1;

architecture behavioral of SEDFFTRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFTRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFTRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFTRX2 : entity is TRUE;
end SEDFFTRX2;

architecture behavioral of SEDFFTRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFTRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFTRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFTRX4 : entity is TRUE;
end SEDFFTRX4;

architecture behavioral of SEDFFTRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFTRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: edff.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity SEDFFTRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_E : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_CK : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_CK : VitalDelayType := DefDummyIsd;
               tisd_E_CK : VitalDelayType := DefDummyIsd;
               ticd_CK : VitalDelayType := DefDummyIcd;
               tpd_CK_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_CK_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tsetup_D_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_E_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_E_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_E_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_E_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_CK : VitalDelayType := DefDummyIsd;
               tsetup_RN_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_RN_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_RN_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SI : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_SE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SI_CK : VitalDelayType := DefDummyIsd;
               tisd_SE_CK : VitalDelayType := DefDummyIsd;
               tsetup_SI_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SI_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SI_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SI_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tsetup_SE_CK_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_SE_CK_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_SE_CK_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_SE_CK_negedge_posedge : VitalDelayType := DefDummyHold;
               tpw_CK_negedge : VitalDelayType := DefDummyWidth;
               tpw_CK_posedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn            : BOOLEAN := DefCombSpikeXOn;
               MsgOn          : BOOLEAN := DefCombSpikeMsgOn;
               instancePath   : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            E : in std_ulogic := 'U';
            SI : in std_ulogic := 'U';
            SE : in std_ulogic := 'U';
            RN : in std_ulogic := 'U'; 
            CK : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of SEDFFTRXL : entity is TRUE;
end SEDFFTRXL;

architecture behavioral of SEDFFTRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL E_dly : std_ulogic := 'X';
     SIGNAL CK_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL SI_dly : std_ulogic := 'X';
     SIGNAL SE_dly : std_ulogic := 'X';

     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL E_ipd : std_ulogic := 'X';
     SIGNAL CK_ipd : std_ulogic := 'X';
     SIGNAL SI_ipd : std_ulogic := 'X';
     SIGNAL SE_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( E_ipd, E, tipd_E );
          VitalWireDelay( CK_ipd, CK, tipd_CK );
          VitalWireDelay( SI_ipd, SI, tipd_SI );
          VitalWireDelay( SE_ipd, SE, tipd_SE );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_CK );
          VitalSignalDelay( E_dly, E_ipd, tisd_E_CK );
          VitalSignalDelay( CK_dly, CK_ipd, ticd_CK );
          VitalSignalDelay( SI_dly, SI_ipd, tisd_SI_CK );
          VitalSignalDelay( SE_dly, SE_ipd, tisd_SE_CK );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_CK );
END BLOCK;

VITALBehavior : PROCESS (D_dly, SI_dly, SE_dly, CK_dly, RN_dly, E_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_CK : std_ulogic := '0';
     VARIABLE TimeMarker_D_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_E_CK : std_ulogic := '0';
     VARIABLE TimeMarker_E_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_CK : std_ulogic := '0';
     VARIABLE TimeMarker_RN_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SI_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SI_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_SE_CK : std_ulogic := '0';
     VARIABLE TimeMarker_SE_CK : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_CK : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_CK : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE S : std_ulogic;
     VARIABLE RNx_dly : std_ulogic := '1';
     VARIABLE SNx_dly : std_ulogic := '1';
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_sedfft_n0 : std_logic_vector( 0 TO 7 );
     VARIABLE n1 : std_ulogic;
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE SEb : std_ulogic;
     VARIABLE scan : std_ulogic;
     VARIABLE flag : std_ulogic;
     VARIABLE Dcheck : std_ulogic;
     VARIABLE DxorSI : std_ulogic;
     VARIABLE Echeck : std_ulogic;
     VARIABLE NoSetReset : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_D_CK_posedge_posedge,
                   SetupLow       => tsetup_D_CK_negedge_posedge,
                   HoldHigh       => thold_D_CK_negedge_posedge,
                   HoldLow        => thold_D_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Dcheck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   TimingData     => TimeMarker_D_CK,
                   Violation      => Tviol_D_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => E_dly,
                   TestSignalName => "E",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_E_CK_posedge_posedge,
                   SetupLow       => tsetup_E_CK_negedge_posedge,
                   HoldHigh       => thold_E_CK_negedge_posedge,
                   HoldLow        => thold_E_CK_posedge_posedge,
                   CheckEnabled   => To_X01(Echeck) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   TimingData     => TimeMarker_E_CK,
                   Violation      => Tviol_E_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SI_dly,
                   TestSignalName => "SI",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SI_CK_posedge_posedge,
                   SetupLow       => tsetup_SI_CK_negedge_posedge,
                   HoldHigh       => thold_SI_CK_negedge_posedge,
                   HoldLow        => thold_SI_CK_posedge_posedge,
                   CheckEnabled   => To_X01(scan) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   TimingData     => TimeMarker_SI_CK,
                   Violation      => Tviol_SI_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SE_dly,
                   TestSignalName => "SE",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_SE_CK_posedge_posedge,
                   SetupLow       => tsetup_SE_CK_negedge_posedge,
                   HoldHigh       => thold_SE_CK_negedge_posedge,
                   HoldLow        => thold_SE_CK_posedge_posedge,
                   CheckEnabled   => To_X01(flag) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   TimingData     => TimeMarker_SE_CK,
                   Violation      => Tviol_SE_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => CK_dly,
                   RefSignalName  => "CK",
                   SetupHigh      => tsetup_RN_CK_posedge_posedge,
                   SetupLow       => tsetup_RN_CK_negedge_posedge,
                   HoldHigh       => thold_RN_CK_negedge_posedge,
                   HoldLow        => thold_RN_CK_posedge_posedge,
                   CheckEnabled   => ((To_X01(SEb) /= '0') and ((To_X01(E_dly) /= '1') or ((To_X01(E_dly) /= '0') and (To_X01(D_dly) /= '0')))),
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   TimingData     => TimeMarker_RN_CK,
                   Violation      => Tviol_RN_CK,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => CK_dly,
                   TestSignalName => "CK",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_CK_posedge,
                   PulseWidthLow  => tpw_CK_negedge,
                   PeriodData     => PeriodCheckInfo_CK,
                   Violation      => PWviol_CK,
                   HeaderMsg      => InstancePath & "/SEDFFTRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := ( 
                       Tviol_D_CK OR 
                       Tviol_RN_CK OR 
                       Tviol_SI_CK OR 
                       Tviol_SE_CK OR 
                       PWviol_CK OR 
                       Tviol_E_CK );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          VitalStateTable ( StateTable => udp_sedfft,
                           DataIn => (NOTIFIER,D_dly,CK_dly,RNx_dly,SNx_dly,E_dly,SI_dly,SE_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_sedfft_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUF( n0 );

          QN_zd := VitalINV( n0 );

          SEb := VitalINV( SE_dly );

          scan := VitalAND3( SE_dly, RNx_dly, SNx_dly );
 
          DxorSI := VitalXOR2(D_dly, SI_dly);

          Dcheck := VitalAND4(SEb,RNx_dly,SNx_dly,E_dly);

          Echeck := VitalAND3(SEb,RNx_dly,SNx_dly);

          flag := VitalAND3(DxorSI,RNx_dly,SNx_dly);

          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_Q,
                             TRUE
                           )
                        ),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( CK_dly'LAST_EVENT,
                             tpd_CK_QN,
                             TRUE
                           )
                        ),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX12 : entity is TRUE;
end TBUFX12;

architecture behavioral of TBUFX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX16 : entity is TRUE;
end TBUFX16;

architecture behavioral of TBUFX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX1 : entity is TRUE;
end TBUFX1;

architecture behavioral of TBUFX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX20 : entity is TRUE;
end TBUFX20;

architecture behavioral of TBUFX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX2 : entity is TRUE;
end TBUFX2;

architecture behavioral of TBUFX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX3 : entity is TRUE;
end TBUFX3;

architecture behavioral of TBUFX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX4 : entity is TRUE;
end TBUFX4;

architecture behavioral of TBUFX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFX8 : entity is TRUE;
end TBUFX8;

architecture behavioral of TBUFX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFXL : entity is TRUE;
end TBUFXL;

architecture behavioral of TBUFXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalBUFIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX12 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX12 : entity is TRUE;
end TBUFIX12;

architecture behavioral of TBUFIX12 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX16 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX16 : entity is TRUE;
end TBUFIX16;

architecture behavioral of TBUFIX16 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX1 : entity is TRUE;
end TBUFIX1;

architecture behavioral of TBUFIX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX20 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX20 : entity is TRUE;
end TBUFIX20;

architecture behavioral of TBUFIX20 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX2 : entity is TRUE;
end TBUFIX2;

architecture behavioral of TBUFIX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX3 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX3 : entity is TRUE;
end TBUFIX3;

architecture behavioral of TBUFIX3 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX4 : entity is TRUE;
end TBUFIX4;

architecture behavioral of TBUFIX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIX8 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIX8 : entity is TRUE;
end TBUFIX8;

architecture behavioral of TBUFIX8 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: inv.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TBUFIXL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_OE_Y : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay)
              );

     port ( 
            OE : in std_ulogic := 'U';
            Y : out std_ulogic;
            A : in std_ulogic := 'U'
           );

     attribute VITAL_LEVEL0 of TBUFIXL : entity is TRUE;
end TBUFIXL;

architecture behavioral of TBUFIXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, OE_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalINVIF1(A_ipd, OE_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_A_Y),
                             TRUE 
                            ),
                      1 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Y),
                             TRUE 
                            )),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tie.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;

entity TIEHI is
 
     port ( Y : out std_ulogic );

     attribute VITAL_LEVEL0 of TIEHI : entity is TRUE;
end TIEHI;

architecture behavioral of TIEHI is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

	signal HIGH : std_ulogic := '1';

BEGIN

-- no timing check section  

-- functionality section 
   VITALBUF (Y, HIGH);

-- no path delay section

end behavioral;
--$Id: tie.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;

entity TIELO is
 
     port ( Y : out std_ulogic );

     attribute VITAL_LEVEL0 of TIELO : entity is TRUE;
end TIELO;

architecture behavioral of TIELO is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;

	signal LOW : std_ulogic := '0';

BEGIN

-- no timing check section  

-- functionality section 
   VITALBUF (Y, LOW);

-- no path delay section

end behavioral;
--$Id: ttlat.genpp,v 1.3 2002/02/13 17:50:55 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TTLATX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_OE_Q : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            OE : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TTLATX1 : entity is TRUE;
end TTLATX1;

architecture behavioral of TTLATX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, OE_ipd, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE xRN_dly : std_ulogic;
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TTLATX1",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TTLATX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          xRN_dly := '1';

          xSN_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUFIF1( n0, OE_ipd );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          SandRandCLK := VitalAND3(xSN_dly,xRN_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_G_Q),
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_D_Q),
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Q),
                             TRUE
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: ttlat.genpp,v 1.3 2002/02/13 17:50:55 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TTLATX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_OE_Q : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            OE : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TTLATX2 : entity is TRUE;
end TTLATX2;

architecture behavioral of TTLATX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, OE_ipd, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE xRN_dly : std_ulogic;
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TTLATX2",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TTLATX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          xRN_dly := '1';

          xSN_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUFIF1( n0, OE_ipd );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          SandRandCLK := VitalAND3(xSN_dly,xRN_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_G_Q),
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_D_Q),
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Q),
                             TRUE
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: ttlat.genpp,v 1.3 2002/02/13 17:50:55 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TTLATX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_OE_Q : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            OE : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TTLATX4 : entity is TRUE;
end TTLATX4;

architecture behavioral of TTLATX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, OE_ipd, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE xRN_dly : std_ulogic;
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TTLATX4",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TTLATX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          xRN_dly := '1';

          xSN_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUFIF1( n0, OE_ipd );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          SandRandCLK := VitalAND3(xSN_dly,xRN_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_G_Q),
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_D_Q),
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Q),
                             TRUE
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: ttlat.genpp,v 1.3 2002/02/13 17:50:55 pearl Exp pearl $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TTLATXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_OE : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_OE_Q : VitalDelayType01Z := (DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay, DefDummyDelay);
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            D : in std_ulogic := 'U';
            OE : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TTLATXL : entity is TRUE;
end TTLATXL;

architecture behavioral of TTLATXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL OE_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( OE_ipd, OE, tipd_OE );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, OE_ipd, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE xRN_dly : std_ulogic;
     VARIABLE xSN_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TTLATXL",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TTLATXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          xRN_dly := '1';

          xSN_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,xRN_dly,xSN_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          Q_zd := VitalBUFIF1( n0, OE_ipd );

          SandR := VitalAND2(xSN_dly,xRN_dly);

          SandRandCLK := VitalAND3(xSN_dly,xRN_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01Z(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_G_Q),
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_D_Q),
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( OE_ipd'LAST_EVENT,
                             VitalExtendToFillDelay(tpd_OE_Q),
                             TRUE
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATX1 : entity is TRUE;
end TLATX1;

architecture behavioral of TLATX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATX1",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATX2 : entity is TRUE;
end TLATX2;

architecture behavioral of TLATX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATX2",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATX4 : entity is TRUE;
end TLATX4;

architecture behavioral of TLATX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATX4",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATXL : entity is TRUE;
end TLATXL;

architecture behavioral of TLATXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATXL",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNX1 : entity is TRUE;
end TLATNX1;

architecture behavioral of TLATNX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNX1",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNX2 : entity is TRUE;
end TLATNX2;

architecture behavioral of TLATNX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNX2",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNX4 : entity is TRUE;
end TLATNX4;

architecture behavioral of TLATNX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNX4",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNXL : entity is TRUE;
end TLATNXL;

architecture behavioral of TLATNXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly)

     -- timing checks section variables
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNXL",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNRX1 : entity is TRUE;
end TLATNRX1;

architecture behavioral of TLATNRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX1",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX1",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNRX2 : entity is TRUE;
end TLATNRX2;

architecture behavioral of TLATNRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX2",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX2",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNRX4 : entity is TRUE;
end TLATNRX4;

architecture behavioral of TLATNRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX4",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRX4",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNRXL : entity is TRUE;
end TLATNRXL;

architecture behavioral of TLATNRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRXL",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNRXL",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSX1 : entity is TRUE;
end TLATNSX1;

architecture behavioral of TLATNSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX1",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX1",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSX2 : entity is TRUE;
end TLATNSX2;

architecture behavioral of TLATNSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX2",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX2",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSX4 : entity is TRUE;
end TLATNSX4;

architecture behavioral of TLATNSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX4",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSX4",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSXL : entity is TRUE;
end TLATNSXL;

architecture behavioral of TLATNSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSXL",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSXL",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSRX1 : entity is TRUE;
end TLATNSRX1;

architecture behavioral of TLATNSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSRX2 : entity is TRUE;
end TLATNSRX2;

architecture behavioral of TLATNSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSRX4 : entity is TRUE;
end TLATNSRX4;

architecture behavioral of TLATNSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATNSRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_GN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_GN : VitalDelayType := DefDummyIsd;
               ticd_GN : VitalDelayType := DefDummyIcd;
               tpd_GN_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_GN_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_GN_negedge : VitalDelayType := DefDummyWidth;
               tsetup_D_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               tsetup_D_GN_negedge_posedge : VitalDelayType := DefDummySetup;
               thold_D_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               thold_D_GN_negedge_posedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_GN : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_RN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_GN : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_GN_posedge_posedge : VitalDelayType := DefDummySetup;
               thold_SN_GN_posedge_posedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            GN : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATNSRXL : entity is TRUE;
end TLATNSRXL;

architecture behavioral of TLATNSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL GN_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL GN_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( GN_ipd, GN, tipd_GN );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_GN );
          VitalSignalDelay( GN_dly, GN_ipd, ticd_GN );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_GN );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_GN );
END BLOCK;

VITALBehavior : PROCESS (D_dly, GN_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_GN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_GN : std_ulogic := '0';
     VARIABLE TimeMarker_D_GN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_GN : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_GN : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_RN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   TimingData     => TimeMarker_RN_GN,
                   Violation      => Tviol_RN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_SN_GN_posedge_posedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_GN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   TimingData     => TimeMarker_SN_GN,
                   Violation      => Tviol_SN_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => GN_dly,
                   RefSignalName  => "GN",
                   SetupHigh      => tsetup_D_GN_posedge_posedge,
                   SetupLow       => tsetup_D_GN_negedge_posedge,
                   HoldHigh       => thold_D_GN_negedge_posedge,
                   HoldLow        => thold_D_GN_posedge_posedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   TimingData     => TimeMarker_D_GN,
                   Violation      => Tviol_D_GN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => GN_dly,
                   TestSignalName => "GN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_GN_negedge,
                   PeriodData     => PeriodCheckInfo_GN,
                   Violation      => PWviol_GN,
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATNSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_GN OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_GN OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_GN OR  
                        PWviol_GN  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalBUF( GN_dly );

          clk := VitalINV( GN_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( GN_dly'LAST_EVENT,
                             tpd_GN_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATRX1 : entity is TRUE;
end TLATRX1;

architecture behavioral of TLATRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX1",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX1",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATRX2 : entity is TRUE;
end TLATRX2;

architecture behavioral of TLATRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX2",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX2",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATRX4 : entity is TRUE;
end TLATRX4;

architecture behavioral of TLATRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX4",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRX4",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATRXL : entity is TRUE;
end TLATRXL;

architecture behavioral of TLATRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRXL",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATRXL",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := '1';

          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSX1 : entity is TRUE;
end TLATSX1;

architecture behavioral of TLATSX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX1",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX1",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSX2 : entity is TRUE;
end TLATSX2;

architecture behavioral of TLATSX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX2",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX2",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSX4 : entity is TRUE;
end TLATSX4;

architecture behavioral of TLATSX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX4",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSX4",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSXL : entity is TRUE;
end TLATSXL;

architecture behavioral of TLATSXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly)

     -- timing checks section variables
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSXL",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSXL",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := '1';

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSRX1 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSRX1 : entity is TRUE;
end TLATSRX1;

architecture behavioral of TLATSRX1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX1",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSRX2 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSRX2 : entity is TRUE;
end TLATSRX2;

architecture behavioral of TLATSRX2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX2",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSRX4 is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSRX4 : entity is TRUE;
end TLATSRX4;

architecture behavioral of TLATSRX4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRX4",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: tlat.genpp,v 1.4 2001/10/02 17:02:07 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity TLATSRXL is

     generic ( tipd_D : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_G : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_D_G : VitalDelayType := DefDummyIsd;
               ticd_G : VitalDelayType := DefDummyIcd;
               tpd_G_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_Q : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_G_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_D_QN : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpw_G_posedge : VitalDelayType := DefDummyWidth;
               tsetup_D_G_posedge_negedge : VitalDelayType := DefDummySetup;
               tsetup_D_G_negedge_negedge : VitalDelayType := DefDummySetup;
               thold_D_G_posedge_negedge : VitalDelayType := DefDummyHold;
               thold_D_G_negedge_negedge : VitalDelayType := DefDummyHold;
               tipd_RN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_RN_G : VitalDelayType := DefDummyIsd;
               tpd_RN_Q : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tpd_RN_QN : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tsetup_RN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_RN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_RN_negedge : VitalDelayType := DefDummyWidth;
               tipd_SN : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tisd_SN_G : VitalDelayType := DefDummyIsd;
               tpd_SN_Q : VitalDelayType01 := (DefDummyDelay, VitalZeroDelay);
               tpd_SN_QN : VitalDelayType01 := (VitalZeroDelay, DefDummyDelay);
               tsetup_SN_G_posedge_negedge : VitalDelayType := DefDummySetup;
               thold_SN_G_posedge_negedge : VitalDelayType := DefDummyHold;
               tpw_SN_negedge : VitalDelayType := DefDummyWidth;
               thold_RN_SN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               thold_SN_RN_posedge_posedge : VitalDelayType := DefDummyRecoverySR;
               TimingChecksOn : BOOLEAN := false;
               XOn : Boolean := DefCombSpikeXOn;
               MsgOn : Boolean := DefCombSpikeMsgOn;
               instancePath : STRING := "*" );

     port ( Q : out std_ulogic;
            QN : out std_ulogic;
            D : in std_ulogic := 'U';
            SN : in std_ulogic := 'U';
            RN : in std_ulogic := 'U';
            G : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of TLATSRXL : entity is TRUE;
end TLATSRXL;

architecture behavioral of TLATSRXL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL D_dly : std_ulogic := 'X';
     SIGNAL G_dly : std_ulogic := 'X';
     SIGNAL SN_dly : std_ulogic := 'X';
     SIGNAL RN_dly : std_ulogic := 'X';
     SIGNAL D_ipd : std_ulogic := 'X';
     SIGNAL G_ipd : std_ulogic := 'X';
     SIGNAL SN_ipd : std_ulogic := 'X';
     SIGNAL RN_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( D_ipd, D, tipd_D );
          VitalWireDelay( G_ipd, G, tipd_G );
          VitalWireDelay( SN_ipd, SN, tipd_SN );
          VitalWireDelay( RN_ipd, RN, tipd_RN );
END BLOCK;

SIGNALDELAY : BLOCK
BEGIN
          VitalSignalDelay( D_dly, D_ipd, tisd_D_G );
          VitalSignalDelay( G_dly, G_ipd, ticd_G );
          VitalSignalDelay( SN_dly, SN_ipd, tisd_SN_G );
          VitalSignalDelay( RN_dly, RN_ipd, tisd_RN_G );
END BLOCK;

VITALBehavior : PROCESS (D_dly, G_dly, SN_dly, RN_dly)

     -- timing checks section variables
     VARIABLE Tviol_RN_G : std_ulogic := '0';
     VARIABLE TimeMarker_RN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_RN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_RN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_SN_G : std_ulogic := '0';
     VARIABLE TimeMarker_SN_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_SN_negedge : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_SN_negedge : VitalPeriodDataType;
     VARIABLE Tviol_D_G : std_ulogic := '0';
     VARIABLE TimeMarker_D_G : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE PWviol_G : std_ulogic := '0';
     VARIABLE PeriodCheckInfo_G : VitalPeriodDataType;
     VARIABLE Tviol_SN_RN : std_ulogic := '0';
     VARIABLE TimeMarker_SN_RN : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tviol_RN_SN : std_ulogic := '0';
     VARIABLE TimeMarker_RN_SN : VitalTimingDataType := VitalTimingDataInit;


     -- functionality section variables
     VARIABLE RNx_dly : std_ulogic;
     VARIABLE SNx_dly : std_ulogic;
     VARIABLE n0 : std_ulogic;
     VARIABLE n0_vec : std_logic_vector( 1 TO 1 );
     VARIABLE PrevData_udp_tlat_n0 : std_logic_vector( 0 TO 4 );
     VARIABLE Q_zd : std_ulogic;
     VARIABLE QN_zd : std_ulogic;
     VARIABLE clk_int : std_ulogic;
     VARIABLE clk : std_ulogic;
     VARIABLE SandR : std_ulogic;
     VARIABLE SandRandCLK : std_ulogic;
     VARIABLE NOTIFIER : std_ulogic := '0';

     -- path delay section variables
     VARIABLE Q_GlitchData : VitalGlitchDataType;
     VARIABLE QN_GlitchData : VitalGlitchDataType;


     BEGIN
          ---------------------------------------------------
          -- Timing checks section
          ---------------------------------------------------
          IF (TimingChecksOn) THEN

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => SN_dly,
                   RefSignalName  => "SN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_SN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   TimingData     => TimeMarker_RN_SN,
                   Violation      => Tviol_RN_SN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => RN_dly,
                   RefSignalName  => "RN",
                   SetupHigh      => 0 ps,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_RN_posedge_posedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'R',
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   TimingData     => TimeMarker_SN_RN,
                   Violation      => Tviol_SN_RN,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_RN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_RN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   TimingData     => TimeMarker_RN_G,
                   Violation      => Tviol_RN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_SN_G_posedge_negedge,
                   SetupLow       => 0 ps,
                   HoldHigh       => 0 ps,
                   HoldLow        => thold_SN_G_posedge_negedge,
                   CheckEnabled   => TRUE,
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   TimingData     => TimeMarker_SN_G,
                   Violation      => Tviol_SN_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalSetupHoldCheck (
                   TestSignal     => D_dly,
                   TestSignalName => "D",
                   RefSignal      => G_dly,
                   RefSignalName  => "G",
                   SetupHigh      => tsetup_D_G_posedge_negedge,
                   SetupLow       => tsetup_D_G_negedge_negedge,
                   HoldHigh       => thold_D_G_negedge_negedge,
                   HoldLow        => thold_D_G_posedge_negedge,
                   CheckEnabled   => To_X01(SandR) /= '0',
                   RefTransition  => 'F',
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   TimingData     => TimeMarker_D_G,
                   Violation      => Tviol_D_G,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => G_dly,
                   TestSignalName => "G",
                   Period         => 0 ps,
                   PulseWidthHigh => tpw_G_posedge,
                   PulseWidthLow  => 0 ps,
                   PeriodData     => PeriodCheckInfo_G,
                   Violation      => PWviol_G,
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   CheckEnabled   => To_X01(SandR) /= '0',
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => SN_dly,
                   TestSignalName => "SN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_SN_negedge,
                   PeriodData     => PeriodCheckInfo_SN_negedge,
                   Violation      => PWviol_SN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

               VitalPeriodPulseCheck (
                   TestSignal     => RN_dly,
                   TestSignalName => "RN",
                   Period         => 0 ps,
                   PulseWidthHigh => 0 ps,
                   PulseWidthLow  => tpw_RN_negedge,
                   PeriodData     => PeriodCheckInfo_RN_negedge,
                   Violation      => PWviol_RN_negedge,
                   HeaderMsg      => InstancePath & "/TLATSRXL",
                   CheckEnabled   => TRUE,
                   XOn            => DefSeqXOn,
                   MsgOn          => DefSeqMsgOn,
                   MsgSeverity    => WARNING );

          END IF;


          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------
          NOTIFIER := (  
                        Tviol_RN_G OR  
                        PWviol_RN_negedge OR
                        Tviol_SN_G OR  
                        PWviol_SN_negedge OR 
                        Tviol_D_G OR  
                        PWviol_G  
                      );

          RNx_dly := RN_dly;

          SNx_dly := SN_dly;


          clk_int := VitalINV( G_dly );

          clk := VitalBUF( G_dly );

          VitalStateTable ( StateTable => udp_tlat,
                           DataIn => (NOTIFIER,D_dly,clk_int,RNx_dly,SNx_dly),
                        NumStates => 1,
                           Result => n0_vec,
                   PreviousDataIn => PrevData_udp_tlat_n0 );
          n0 := n0_vec(1);

          QN_zd := VitalINV( n0 );

          Q_zd := VitalBUF( n0 );

          SandR := VitalAND2(SNx_dly,RNx_dly);

          SandRandCLK := VitalAND3(SNx_dly,RNx_dly,clk);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Q,
               OutSignalName => "Q",
               OutTemp => Q_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_Q,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_Q,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_Q,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_Q,
                             TRUE 
                           )),
               GlitchData => Q_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

          VitalPathDelay01(
               OutSignal => QN,
               OutSignalName => "QN",
               OutTemp => QN_zd,
               Paths => (
                      0 => ( G_dly'LAST_EVENT,
                             tpd_G_QN,
                             ( To_X01(SandR) ) /= '0' 
                           ),
                      1 => ( D_dly'LAST_EVENT,
                             tpd_D_QN,
                             ( To_X01(SandRandCLK) ) /= '0' 
                           ),
                      2 => ( SN_dly'LAST_EVENT,
                             tpd_SN_QN,
                             TRUE 
                           ),
                      3 => ( RN_dly'LAST_EVENT,
                             tpd_RN_QN,
                             TRUE 
                           )),
               GlitchData => QN_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR2X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR2X1 : entity is TRUE;
end XNOR2X1;

architecture behavioral of XNOR2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR2X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR2X2 : entity is TRUE;
end XNOR2X2;

architecture behavioral of XNOR2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR2X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR2X4 : entity is TRUE;
end XNOR2X4;

architecture behavioral of XNOR2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XNOR2XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XNOR2XL : entity is TRUE;
end XNOR2XL;

architecture behavioral of XNOR2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXNOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR2X1 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR2X1 : entity is TRUE;
end XOR2X1;

architecture behavioral of XOR2X1 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR2X2 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR2X2 : entity is TRUE;
end XOR2X2;

architecture behavioral of XOR2X2 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR2X4 is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR2X4 : entity is TRUE;
end XOR2X4;

architecture behavioral of XOR2X4 is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;
--$Id: xor.genpp,v 1.2 2001/06/25 18:00:42 pearl Exp $
--CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF ARTISAN COMPONENTS, INC.
--
--Copyright (c) 2002 Artisan Components, Inc.  All Rights Reserved.
--
--Use of this Software/Data is subject to the terms and conditions of
--the applicable license agreement between Artisan Components, Inc. and
--TSMC.  In addition, this Software/Data
--is protected by copyright law and international treaties.
--
--The copyright notice(s) in this Software/Data does not indicate actual
--or intended publication of this Software/Data.

LIBRARY IEEE;
USE IEEE.Std_logic_1164.all;
USE IEEE.VITAL_Timing.all;
USE IEEE.VITAL_Primitives.all;
USE work.prim.all;

entity XOR2XL is

     generic ( 
               XOn    : BOOLEAN := DefCombSpikeXOn;
               MsgOn  : BOOLEAN := DefCombSpikeMsgOn;
               InstancePath : STRING := "*";
               tipd_A : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tipd_B : VitalDelayType01 := (DefDummyIpd, DefDummyIpd);
               tpd_A_Y_B_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y_B_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_A_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_0 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y_A_EQ_1 : VitalDelayType01 := (DefDummyDelay, DefDummyDelay);
               tpd_B_Y : VitalDelayType01 := (DefDummyDelay, DefDummyDelay));

     port ( Y : out std_ulogic;
            A : in std_ulogic := 'U';
            B : in std_ulogic := 'U' );

     attribute VITAL_LEVEL0 of XOR2XL : entity is TRUE;
end XOR2XL;

architecture behavioral of XOR2XL is
     attribute VITAL_LEVEL1 of behavioral : architecture is TRUE;


     SIGNAL A_ipd : std_ulogic := 'X';
     SIGNAL B_ipd : std_ulogic := 'X';

BEGIN

---------------------------------------------------
-- Input Path Delays
---------------------------------------------------
WIREDELAY : BLOCK
BEGIN
          VitalWireDelay( A_ipd, A, tipd_A );
          VitalWireDelay( B_ipd, B, tipd_B );
END BLOCK;

VITALBehavior : PROCESS (A_ipd, B_ipd)


     -- functionality section variables
     VARIABLE Y_zd : std_ulogic;

     -- path delay section variables
     VARIABLE Y_GlitchData : VitalGlitchDataType;


     BEGIN

          ---------------------------------------------------
          -- Functionality section
          ---------------------------------------------------

          Y_zd := VitalXOR2(A_ipd,B_ipd);


          ---------------------------------------------------
          -- Path delay section
          ---------------------------------------------------
          VitalPathDelay01(
               OutSignal => Y,
               OutSignalName => "Y",
               OutTemp => Y_zd,
               Paths => (
                      0 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_0,
                             (To_X01(B_ipd) /= '1')),
                      1 => ( A_ipd'LAST_EVENT,
                             tpd_A_Y_B_EQ_1,
                             (To_X01(B_ipd) /= '0')),
                      2 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_0,
                             (To_X01(A_ipd) /= '1')),
                      3 => ( B_ipd'LAST_EVENT,
                             tpd_B_Y_A_EQ_1,
                             (To_X01(A_ipd) /= '0'))),
               GlitchData => Y_GlitchData,
               Mode  => OnEvent,
               XOn => XOn,
               MsgOn => MsgOn,
               MsgSeverity => WARNING);

END PROCESS;
end behavioral;